module  tryfunct2( 
	input 
);
