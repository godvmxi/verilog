//megafunction wizard: %Altera SOPC Builder%
//GENERATION: STANDARD
//VERSION: WM1.0


//Legal Notice: (C)2015 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module PIO_LCD_B_s1_arbitrator (
                                 // inputs:
                                  PIO_LCD_B_s1_readdata,
                                  clk,
                                  cpu_data_master_address_to_slave,
                                  cpu_data_master_read,
                                  cpu_data_master_waitrequest,
                                  cpu_data_master_write,
                                  cpu_data_master_writedata,
                                  reset_n,

                                 // outputs:
                                  PIO_LCD_B_s1_address,
                                  PIO_LCD_B_s1_chipselect,
                                  PIO_LCD_B_s1_readdata_from_sa,
                                  PIO_LCD_B_s1_reset_n,
                                  PIO_LCD_B_s1_write_n,
                                  PIO_LCD_B_s1_writedata,
                                  cpu_data_master_granted_PIO_LCD_B_s1,
                                  cpu_data_master_qualified_request_PIO_LCD_B_s1,
                                  cpu_data_master_read_data_valid_PIO_LCD_B_s1,
                                  cpu_data_master_requests_PIO_LCD_B_s1,
                                  d1_PIO_LCD_B_s1_end_xfer
                               )
;

  output  [  1: 0] PIO_LCD_B_s1_address;
  output           PIO_LCD_B_s1_chipselect;
  output  [ 31: 0] PIO_LCD_B_s1_readdata_from_sa;
  output           PIO_LCD_B_s1_reset_n;
  output           PIO_LCD_B_s1_write_n;
  output  [ 31: 0] PIO_LCD_B_s1_writedata;
  output           cpu_data_master_granted_PIO_LCD_B_s1;
  output           cpu_data_master_qualified_request_PIO_LCD_B_s1;
  output           cpu_data_master_read_data_valid_PIO_LCD_B_s1;
  output           cpu_data_master_requests_PIO_LCD_B_s1;
  output           d1_PIO_LCD_B_s1_end_xfer;
  input   [ 31: 0] PIO_LCD_B_s1_readdata;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_read;
  input            cpu_data_master_waitrequest;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;

  wire    [  1: 0] PIO_LCD_B_s1_address;
  wire             PIO_LCD_B_s1_allgrants;
  wire             PIO_LCD_B_s1_allow_new_arb_cycle;
  wire             PIO_LCD_B_s1_any_bursting_master_saved_grant;
  wire             PIO_LCD_B_s1_any_continuerequest;
  wire             PIO_LCD_B_s1_arb_counter_enable;
  reg     [  1: 0] PIO_LCD_B_s1_arb_share_counter;
  wire    [  1: 0] PIO_LCD_B_s1_arb_share_counter_next_value;
  wire    [  1: 0] PIO_LCD_B_s1_arb_share_set_values;
  wire             PIO_LCD_B_s1_beginbursttransfer_internal;
  wire             PIO_LCD_B_s1_begins_xfer;
  wire             PIO_LCD_B_s1_chipselect;
  wire             PIO_LCD_B_s1_end_xfer;
  wire             PIO_LCD_B_s1_firsttransfer;
  wire             PIO_LCD_B_s1_grant_vector;
  wire             PIO_LCD_B_s1_in_a_read_cycle;
  wire             PIO_LCD_B_s1_in_a_write_cycle;
  wire             PIO_LCD_B_s1_master_qreq_vector;
  wire             PIO_LCD_B_s1_non_bursting_master_requests;
  wire    [ 31: 0] PIO_LCD_B_s1_readdata_from_sa;
  reg              PIO_LCD_B_s1_reg_firsttransfer;
  wire             PIO_LCD_B_s1_reset_n;
  reg              PIO_LCD_B_s1_slavearbiterlockenable;
  wire             PIO_LCD_B_s1_slavearbiterlockenable2;
  wire             PIO_LCD_B_s1_unreg_firsttransfer;
  wire             PIO_LCD_B_s1_waits_for_read;
  wire             PIO_LCD_B_s1_waits_for_write;
  wire             PIO_LCD_B_s1_write_n;
  wire    [ 31: 0] PIO_LCD_B_s1_writedata;
  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_PIO_LCD_B_s1;
  wire             cpu_data_master_qualified_request_PIO_LCD_B_s1;
  wire             cpu_data_master_read_data_valid_PIO_LCD_B_s1;
  wire             cpu_data_master_requests_PIO_LCD_B_s1;
  wire             cpu_data_master_saved_grant_PIO_LCD_B_s1;
  reg              d1_PIO_LCD_B_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_PIO_LCD_B_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 26: 0] shifted_address_to_PIO_LCD_B_s1_from_cpu_data_master;
  wire             wait_for_PIO_LCD_B_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~PIO_LCD_B_s1_end_xfer;
    end


  assign PIO_LCD_B_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_PIO_LCD_B_s1));
  //assign PIO_LCD_B_s1_readdata_from_sa = PIO_LCD_B_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign PIO_LCD_B_s1_readdata_from_sa = PIO_LCD_B_s1_readdata;

  assign cpu_data_master_requests_PIO_LCD_B_s1 = ({cpu_data_master_address_to_slave[26 : 4] , 4'b0} == 27'h1840) & (cpu_data_master_read | cpu_data_master_write);
  //PIO_LCD_B_s1_arb_share_counter set values, which is an e_mux
  assign PIO_LCD_B_s1_arb_share_set_values = 1;

  //PIO_LCD_B_s1_non_bursting_master_requests mux, which is an e_mux
  assign PIO_LCD_B_s1_non_bursting_master_requests = cpu_data_master_requests_PIO_LCD_B_s1;

  //PIO_LCD_B_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign PIO_LCD_B_s1_any_bursting_master_saved_grant = 0;

  //PIO_LCD_B_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign PIO_LCD_B_s1_arb_share_counter_next_value = PIO_LCD_B_s1_firsttransfer ? (PIO_LCD_B_s1_arb_share_set_values - 1) : |PIO_LCD_B_s1_arb_share_counter ? (PIO_LCD_B_s1_arb_share_counter - 1) : 0;

  //PIO_LCD_B_s1_allgrants all slave grants, which is an e_mux
  assign PIO_LCD_B_s1_allgrants = |PIO_LCD_B_s1_grant_vector;

  //PIO_LCD_B_s1_end_xfer assignment, which is an e_assign
  assign PIO_LCD_B_s1_end_xfer = ~(PIO_LCD_B_s1_waits_for_read | PIO_LCD_B_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_PIO_LCD_B_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_PIO_LCD_B_s1 = PIO_LCD_B_s1_end_xfer & (~PIO_LCD_B_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //PIO_LCD_B_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign PIO_LCD_B_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_PIO_LCD_B_s1 & PIO_LCD_B_s1_allgrants) | (end_xfer_arb_share_counter_term_PIO_LCD_B_s1 & ~PIO_LCD_B_s1_non_bursting_master_requests);

  //PIO_LCD_B_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_B_s1_arb_share_counter <= 0;
      else if (PIO_LCD_B_s1_arb_counter_enable)
          PIO_LCD_B_s1_arb_share_counter <= PIO_LCD_B_s1_arb_share_counter_next_value;
    end


  //PIO_LCD_B_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_B_s1_slavearbiterlockenable <= 0;
      else if ((|PIO_LCD_B_s1_master_qreq_vector & end_xfer_arb_share_counter_term_PIO_LCD_B_s1) | (end_xfer_arb_share_counter_term_PIO_LCD_B_s1 & ~PIO_LCD_B_s1_non_bursting_master_requests))
          PIO_LCD_B_s1_slavearbiterlockenable <= |PIO_LCD_B_s1_arb_share_counter_next_value;
    end


  //cpu/data_master PIO_LCD_B/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = PIO_LCD_B_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //PIO_LCD_B_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign PIO_LCD_B_s1_slavearbiterlockenable2 = |PIO_LCD_B_s1_arb_share_counter_next_value;

  //cpu/data_master PIO_LCD_B/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = PIO_LCD_B_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //PIO_LCD_B_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign PIO_LCD_B_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_PIO_LCD_B_s1 = cpu_data_master_requests_PIO_LCD_B_s1 & ~(((~cpu_data_master_waitrequest) & cpu_data_master_write));
  //PIO_LCD_B_s1_writedata mux, which is an e_mux
  assign PIO_LCD_B_s1_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_PIO_LCD_B_s1 = cpu_data_master_qualified_request_PIO_LCD_B_s1;

  //cpu/data_master saved-grant PIO_LCD_B/s1, which is an e_assign
  assign cpu_data_master_saved_grant_PIO_LCD_B_s1 = cpu_data_master_requests_PIO_LCD_B_s1;

  //allow new arb cycle for PIO_LCD_B/s1, which is an e_assign
  assign PIO_LCD_B_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign PIO_LCD_B_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign PIO_LCD_B_s1_master_qreq_vector = 1;

  //PIO_LCD_B_s1_reset_n assignment, which is an e_assign
  assign PIO_LCD_B_s1_reset_n = reset_n;

  assign PIO_LCD_B_s1_chipselect = cpu_data_master_granted_PIO_LCD_B_s1;
  //PIO_LCD_B_s1_firsttransfer first transaction, which is an e_assign
  assign PIO_LCD_B_s1_firsttransfer = PIO_LCD_B_s1_begins_xfer ? PIO_LCD_B_s1_unreg_firsttransfer : PIO_LCD_B_s1_reg_firsttransfer;

  //PIO_LCD_B_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign PIO_LCD_B_s1_unreg_firsttransfer = ~(PIO_LCD_B_s1_slavearbiterlockenable & PIO_LCD_B_s1_any_continuerequest);

  //PIO_LCD_B_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_B_s1_reg_firsttransfer <= 1'b1;
      else if (PIO_LCD_B_s1_begins_xfer)
          PIO_LCD_B_s1_reg_firsttransfer <= PIO_LCD_B_s1_unreg_firsttransfer;
    end


  //PIO_LCD_B_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign PIO_LCD_B_s1_beginbursttransfer_internal = PIO_LCD_B_s1_begins_xfer;

  //~PIO_LCD_B_s1_write_n assignment, which is an e_mux
  assign PIO_LCD_B_s1_write_n = ~(cpu_data_master_granted_PIO_LCD_B_s1 & cpu_data_master_write);

  assign shifted_address_to_PIO_LCD_B_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //PIO_LCD_B_s1_address mux, which is an e_mux
  assign PIO_LCD_B_s1_address = shifted_address_to_PIO_LCD_B_s1_from_cpu_data_master >> 2;

  //d1_PIO_LCD_B_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_PIO_LCD_B_s1_end_xfer <= 1;
      else 
        d1_PIO_LCD_B_s1_end_xfer <= PIO_LCD_B_s1_end_xfer;
    end


  //PIO_LCD_B_s1_waits_for_read in a cycle, which is an e_mux
  assign PIO_LCD_B_s1_waits_for_read = PIO_LCD_B_s1_in_a_read_cycle & PIO_LCD_B_s1_begins_xfer;

  //PIO_LCD_B_s1_in_a_read_cycle assignment, which is an e_assign
  assign PIO_LCD_B_s1_in_a_read_cycle = cpu_data_master_granted_PIO_LCD_B_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = PIO_LCD_B_s1_in_a_read_cycle;

  //PIO_LCD_B_s1_waits_for_write in a cycle, which is an e_mux
  assign PIO_LCD_B_s1_waits_for_write = PIO_LCD_B_s1_in_a_write_cycle & 0;

  //PIO_LCD_B_s1_in_a_write_cycle assignment, which is an e_assign
  assign PIO_LCD_B_s1_in_a_write_cycle = cpu_data_master_granted_PIO_LCD_B_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = PIO_LCD_B_s1_in_a_write_cycle;

  assign wait_for_PIO_LCD_B_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //PIO_LCD_B/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module PIO_LCD_CLK_s1_arbitrator (
                                   // inputs:
                                    PIO_LCD_CLK_s1_readdata,
                                    clk,
                                    cpu_data_master_address_to_slave,
                                    cpu_data_master_read,
                                    cpu_data_master_waitrequest,
                                    cpu_data_master_write,
                                    cpu_data_master_writedata,
                                    reset_n,

                                   // outputs:
                                    PIO_LCD_CLK_s1_address,
                                    PIO_LCD_CLK_s1_chipselect,
                                    PIO_LCD_CLK_s1_readdata_from_sa,
                                    PIO_LCD_CLK_s1_reset_n,
                                    PIO_LCD_CLK_s1_write_n,
                                    PIO_LCD_CLK_s1_writedata,
                                    cpu_data_master_granted_PIO_LCD_CLK_s1,
                                    cpu_data_master_qualified_request_PIO_LCD_CLK_s1,
                                    cpu_data_master_read_data_valid_PIO_LCD_CLK_s1,
                                    cpu_data_master_requests_PIO_LCD_CLK_s1,
                                    d1_PIO_LCD_CLK_s1_end_xfer
                                 )
;

  output  [  1: 0] PIO_LCD_CLK_s1_address;
  output           PIO_LCD_CLK_s1_chipselect;
  output  [ 31: 0] PIO_LCD_CLK_s1_readdata_from_sa;
  output           PIO_LCD_CLK_s1_reset_n;
  output           PIO_LCD_CLK_s1_write_n;
  output  [ 31: 0] PIO_LCD_CLK_s1_writedata;
  output           cpu_data_master_granted_PIO_LCD_CLK_s1;
  output           cpu_data_master_qualified_request_PIO_LCD_CLK_s1;
  output           cpu_data_master_read_data_valid_PIO_LCD_CLK_s1;
  output           cpu_data_master_requests_PIO_LCD_CLK_s1;
  output           d1_PIO_LCD_CLK_s1_end_xfer;
  input   [ 31: 0] PIO_LCD_CLK_s1_readdata;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_read;
  input            cpu_data_master_waitrequest;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;

  wire    [  1: 0] PIO_LCD_CLK_s1_address;
  wire             PIO_LCD_CLK_s1_allgrants;
  wire             PIO_LCD_CLK_s1_allow_new_arb_cycle;
  wire             PIO_LCD_CLK_s1_any_bursting_master_saved_grant;
  wire             PIO_LCD_CLK_s1_any_continuerequest;
  wire             PIO_LCD_CLK_s1_arb_counter_enable;
  reg     [  1: 0] PIO_LCD_CLK_s1_arb_share_counter;
  wire    [  1: 0] PIO_LCD_CLK_s1_arb_share_counter_next_value;
  wire    [  1: 0] PIO_LCD_CLK_s1_arb_share_set_values;
  wire             PIO_LCD_CLK_s1_beginbursttransfer_internal;
  wire             PIO_LCD_CLK_s1_begins_xfer;
  wire             PIO_LCD_CLK_s1_chipselect;
  wire             PIO_LCD_CLK_s1_end_xfer;
  wire             PIO_LCD_CLK_s1_firsttransfer;
  wire             PIO_LCD_CLK_s1_grant_vector;
  wire             PIO_LCD_CLK_s1_in_a_read_cycle;
  wire             PIO_LCD_CLK_s1_in_a_write_cycle;
  wire             PIO_LCD_CLK_s1_master_qreq_vector;
  wire             PIO_LCD_CLK_s1_non_bursting_master_requests;
  wire    [ 31: 0] PIO_LCD_CLK_s1_readdata_from_sa;
  reg              PIO_LCD_CLK_s1_reg_firsttransfer;
  wire             PIO_LCD_CLK_s1_reset_n;
  reg              PIO_LCD_CLK_s1_slavearbiterlockenable;
  wire             PIO_LCD_CLK_s1_slavearbiterlockenable2;
  wire             PIO_LCD_CLK_s1_unreg_firsttransfer;
  wire             PIO_LCD_CLK_s1_waits_for_read;
  wire             PIO_LCD_CLK_s1_waits_for_write;
  wire             PIO_LCD_CLK_s1_write_n;
  wire    [ 31: 0] PIO_LCD_CLK_s1_writedata;
  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_PIO_LCD_CLK_s1;
  wire             cpu_data_master_qualified_request_PIO_LCD_CLK_s1;
  wire             cpu_data_master_read_data_valid_PIO_LCD_CLK_s1;
  wire             cpu_data_master_requests_PIO_LCD_CLK_s1;
  wire             cpu_data_master_saved_grant_PIO_LCD_CLK_s1;
  reg              d1_PIO_LCD_CLK_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_PIO_LCD_CLK_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 26: 0] shifted_address_to_PIO_LCD_CLK_s1_from_cpu_data_master;
  wire             wait_for_PIO_LCD_CLK_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~PIO_LCD_CLK_s1_end_xfer;
    end


  assign PIO_LCD_CLK_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_PIO_LCD_CLK_s1));
  //assign PIO_LCD_CLK_s1_readdata_from_sa = PIO_LCD_CLK_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign PIO_LCD_CLK_s1_readdata_from_sa = PIO_LCD_CLK_s1_readdata;

  assign cpu_data_master_requests_PIO_LCD_CLK_s1 = ({cpu_data_master_address_to_slave[26 : 4] , 4'b0} == 27'h1870) & (cpu_data_master_read | cpu_data_master_write);
  //PIO_LCD_CLK_s1_arb_share_counter set values, which is an e_mux
  assign PIO_LCD_CLK_s1_arb_share_set_values = 1;

  //PIO_LCD_CLK_s1_non_bursting_master_requests mux, which is an e_mux
  assign PIO_LCD_CLK_s1_non_bursting_master_requests = cpu_data_master_requests_PIO_LCD_CLK_s1;

  //PIO_LCD_CLK_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign PIO_LCD_CLK_s1_any_bursting_master_saved_grant = 0;

  //PIO_LCD_CLK_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign PIO_LCD_CLK_s1_arb_share_counter_next_value = PIO_LCD_CLK_s1_firsttransfer ? (PIO_LCD_CLK_s1_arb_share_set_values - 1) : |PIO_LCD_CLK_s1_arb_share_counter ? (PIO_LCD_CLK_s1_arb_share_counter - 1) : 0;

  //PIO_LCD_CLK_s1_allgrants all slave grants, which is an e_mux
  assign PIO_LCD_CLK_s1_allgrants = |PIO_LCD_CLK_s1_grant_vector;

  //PIO_LCD_CLK_s1_end_xfer assignment, which is an e_assign
  assign PIO_LCD_CLK_s1_end_xfer = ~(PIO_LCD_CLK_s1_waits_for_read | PIO_LCD_CLK_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_PIO_LCD_CLK_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_PIO_LCD_CLK_s1 = PIO_LCD_CLK_s1_end_xfer & (~PIO_LCD_CLK_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //PIO_LCD_CLK_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign PIO_LCD_CLK_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_PIO_LCD_CLK_s1 & PIO_LCD_CLK_s1_allgrants) | (end_xfer_arb_share_counter_term_PIO_LCD_CLK_s1 & ~PIO_LCD_CLK_s1_non_bursting_master_requests);

  //PIO_LCD_CLK_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_CLK_s1_arb_share_counter <= 0;
      else if (PIO_LCD_CLK_s1_arb_counter_enable)
          PIO_LCD_CLK_s1_arb_share_counter <= PIO_LCD_CLK_s1_arb_share_counter_next_value;
    end


  //PIO_LCD_CLK_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_CLK_s1_slavearbiterlockenable <= 0;
      else if ((|PIO_LCD_CLK_s1_master_qreq_vector & end_xfer_arb_share_counter_term_PIO_LCD_CLK_s1) | (end_xfer_arb_share_counter_term_PIO_LCD_CLK_s1 & ~PIO_LCD_CLK_s1_non_bursting_master_requests))
          PIO_LCD_CLK_s1_slavearbiterlockenable <= |PIO_LCD_CLK_s1_arb_share_counter_next_value;
    end


  //cpu/data_master PIO_LCD_CLK/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = PIO_LCD_CLK_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //PIO_LCD_CLK_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign PIO_LCD_CLK_s1_slavearbiterlockenable2 = |PIO_LCD_CLK_s1_arb_share_counter_next_value;

  //cpu/data_master PIO_LCD_CLK/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = PIO_LCD_CLK_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //PIO_LCD_CLK_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign PIO_LCD_CLK_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_PIO_LCD_CLK_s1 = cpu_data_master_requests_PIO_LCD_CLK_s1 & ~(((~cpu_data_master_waitrequest) & cpu_data_master_write));
  //PIO_LCD_CLK_s1_writedata mux, which is an e_mux
  assign PIO_LCD_CLK_s1_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_PIO_LCD_CLK_s1 = cpu_data_master_qualified_request_PIO_LCD_CLK_s1;

  //cpu/data_master saved-grant PIO_LCD_CLK/s1, which is an e_assign
  assign cpu_data_master_saved_grant_PIO_LCD_CLK_s1 = cpu_data_master_requests_PIO_LCD_CLK_s1;

  //allow new arb cycle for PIO_LCD_CLK/s1, which is an e_assign
  assign PIO_LCD_CLK_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign PIO_LCD_CLK_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign PIO_LCD_CLK_s1_master_qreq_vector = 1;

  //PIO_LCD_CLK_s1_reset_n assignment, which is an e_assign
  assign PIO_LCD_CLK_s1_reset_n = reset_n;

  assign PIO_LCD_CLK_s1_chipselect = cpu_data_master_granted_PIO_LCD_CLK_s1;
  //PIO_LCD_CLK_s1_firsttransfer first transaction, which is an e_assign
  assign PIO_LCD_CLK_s1_firsttransfer = PIO_LCD_CLK_s1_begins_xfer ? PIO_LCD_CLK_s1_unreg_firsttransfer : PIO_LCD_CLK_s1_reg_firsttransfer;

  //PIO_LCD_CLK_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign PIO_LCD_CLK_s1_unreg_firsttransfer = ~(PIO_LCD_CLK_s1_slavearbiterlockenable & PIO_LCD_CLK_s1_any_continuerequest);

  //PIO_LCD_CLK_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_CLK_s1_reg_firsttransfer <= 1'b1;
      else if (PIO_LCD_CLK_s1_begins_xfer)
          PIO_LCD_CLK_s1_reg_firsttransfer <= PIO_LCD_CLK_s1_unreg_firsttransfer;
    end


  //PIO_LCD_CLK_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign PIO_LCD_CLK_s1_beginbursttransfer_internal = PIO_LCD_CLK_s1_begins_xfer;

  //~PIO_LCD_CLK_s1_write_n assignment, which is an e_mux
  assign PIO_LCD_CLK_s1_write_n = ~(cpu_data_master_granted_PIO_LCD_CLK_s1 & cpu_data_master_write);

  assign shifted_address_to_PIO_LCD_CLK_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //PIO_LCD_CLK_s1_address mux, which is an e_mux
  assign PIO_LCD_CLK_s1_address = shifted_address_to_PIO_LCD_CLK_s1_from_cpu_data_master >> 2;

  //d1_PIO_LCD_CLK_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_PIO_LCD_CLK_s1_end_xfer <= 1;
      else 
        d1_PIO_LCD_CLK_s1_end_xfer <= PIO_LCD_CLK_s1_end_xfer;
    end


  //PIO_LCD_CLK_s1_waits_for_read in a cycle, which is an e_mux
  assign PIO_LCD_CLK_s1_waits_for_read = PIO_LCD_CLK_s1_in_a_read_cycle & PIO_LCD_CLK_s1_begins_xfer;

  //PIO_LCD_CLK_s1_in_a_read_cycle assignment, which is an e_assign
  assign PIO_LCD_CLK_s1_in_a_read_cycle = cpu_data_master_granted_PIO_LCD_CLK_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = PIO_LCD_CLK_s1_in_a_read_cycle;

  //PIO_LCD_CLK_s1_waits_for_write in a cycle, which is an e_mux
  assign PIO_LCD_CLK_s1_waits_for_write = PIO_LCD_CLK_s1_in_a_write_cycle & 0;

  //PIO_LCD_CLK_s1_in_a_write_cycle assignment, which is an e_assign
  assign PIO_LCD_CLK_s1_in_a_write_cycle = cpu_data_master_granted_PIO_LCD_CLK_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = PIO_LCD_CLK_s1_in_a_write_cycle;

  assign wait_for_PIO_LCD_CLK_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //PIO_LCD_CLK/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module PIO_LCD_CTRL_s1_arbitrator (
                                    // inputs:
                                     PIO_LCD_CTRL_s1_readdata,
                                     clk,
                                     cpu_data_master_address_to_slave,
                                     cpu_data_master_read,
                                     cpu_data_master_waitrequest,
                                     cpu_data_master_write,
                                     cpu_data_master_writedata,
                                     reset_n,

                                    // outputs:
                                     PIO_LCD_CTRL_s1_address,
                                     PIO_LCD_CTRL_s1_chipselect,
                                     PIO_LCD_CTRL_s1_readdata_from_sa,
                                     PIO_LCD_CTRL_s1_reset_n,
                                     PIO_LCD_CTRL_s1_write_n,
                                     PIO_LCD_CTRL_s1_writedata,
                                     cpu_data_master_granted_PIO_LCD_CTRL_s1,
                                     cpu_data_master_qualified_request_PIO_LCD_CTRL_s1,
                                     cpu_data_master_read_data_valid_PIO_LCD_CTRL_s1,
                                     cpu_data_master_requests_PIO_LCD_CTRL_s1,
                                     d1_PIO_LCD_CTRL_s1_end_xfer
                                  )
;

  output  [  1: 0] PIO_LCD_CTRL_s1_address;
  output           PIO_LCD_CTRL_s1_chipselect;
  output  [ 31: 0] PIO_LCD_CTRL_s1_readdata_from_sa;
  output           PIO_LCD_CTRL_s1_reset_n;
  output           PIO_LCD_CTRL_s1_write_n;
  output  [ 31: 0] PIO_LCD_CTRL_s1_writedata;
  output           cpu_data_master_granted_PIO_LCD_CTRL_s1;
  output           cpu_data_master_qualified_request_PIO_LCD_CTRL_s1;
  output           cpu_data_master_read_data_valid_PIO_LCD_CTRL_s1;
  output           cpu_data_master_requests_PIO_LCD_CTRL_s1;
  output           d1_PIO_LCD_CTRL_s1_end_xfer;
  input   [ 31: 0] PIO_LCD_CTRL_s1_readdata;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_read;
  input            cpu_data_master_waitrequest;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;

  wire    [  1: 0] PIO_LCD_CTRL_s1_address;
  wire             PIO_LCD_CTRL_s1_allgrants;
  wire             PIO_LCD_CTRL_s1_allow_new_arb_cycle;
  wire             PIO_LCD_CTRL_s1_any_bursting_master_saved_grant;
  wire             PIO_LCD_CTRL_s1_any_continuerequest;
  wire             PIO_LCD_CTRL_s1_arb_counter_enable;
  reg     [  1: 0] PIO_LCD_CTRL_s1_arb_share_counter;
  wire    [  1: 0] PIO_LCD_CTRL_s1_arb_share_counter_next_value;
  wire    [  1: 0] PIO_LCD_CTRL_s1_arb_share_set_values;
  wire             PIO_LCD_CTRL_s1_beginbursttransfer_internal;
  wire             PIO_LCD_CTRL_s1_begins_xfer;
  wire             PIO_LCD_CTRL_s1_chipselect;
  wire             PIO_LCD_CTRL_s1_end_xfer;
  wire             PIO_LCD_CTRL_s1_firsttransfer;
  wire             PIO_LCD_CTRL_s1_grant_vector;
  wire             PIO_LCD_CTRL_s1_in_a_read_cycle;
  wire             PIO_LCD_CTRL_s1_in_a_write_cycle;
  wire             PIO_LCD_CTRL_s1_master_qreq_vector;
  wire             PIO_LCD_CTRL_s1_non_bursting_master_requests;
  wire    [ 31: 0] PIO_LCD_CTRL_s1_readdata_from_sa;
  reg              PIO_LCD_CTRL_s1_reg_firsttransfer;
  wire             PIO_LCD_CTRL_s1_reset_n;
  reg              PIO_LCD_CTRL_s1_slavearbiterlockenable;
  wire             PIO_LCD_CTRL_s1_slavearbiterlockenable2;
  wire             PIO_LCD_CTRL_s1_unreg_firsttransfer;
  wire             PIO_LCD_CTRL_s1_waits_for_read;
  wire             PIO_LCD_CTRL_s1_waits_for_write;
  wire             PIO_LCD_CTRL_s1_write_n;
  wire    [ 31: 0] PIO_LCD_CTRL_s1_writedata;
  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_PIO_LCD_CTRL_s1;
  wire             cpu_data_master_qualified_request_PIO_LCD_CTRL_s1;
  wire             cpu_data_master_read_data_valid_PIO_LCD_CTRL_s1;
  wire             cpu_data_master_requests_PIO_LCD_CTRL_s1;
  wire             cpu_data_master_saved_grant_PIO_LCD_CTRL_s1;
  reg              d1_PIO_LCD_CTRL_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_PIO_LCD_CTRL_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 26: 0] shifted_address_to_PIO_LCD_CTRL_s1_from_cpu_data_master;
  wire             wait_for_PIO_LCD_CTRL_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~PIO_LCD_CTRL_s1_end_xfer;
    end


  assign PIO_LCD_CTRL_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_PIO_LCD_CTRL_s1));
  //assign PIO_LCD_CTRL_s1_readdata_from_sa = PIO_LCD_CTRL_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign PIO_LCD_CTRL_s1_readdata_from_sa = PIO_LCD_CTRL_s1_readdata;

  assign cpu_data_master_requests_PIO_LCD_CTRL_s1 = ({cpu_data_master_address_to_slave[26 : 4] , 4'b0} == 27'h1830) & (cpu_data_master_read | cpu_data_master_write);
  //PIO_LCD_CTRL_s1_arb_share_counter set values, which is an e_mux
  assign PIO_LCD_CTRL_s1_arb_share_set_values = 1;

  //PIO_LCD_CTRL_s1_non_bursting_master_requests mux, which is an e_mux
  assign PIO_LCD_CTRL_s1_non_bursting_master_requests = cpu_data_master_requests_PIO_LCD_CTRL_s1;

  //PIO_LCD_CTRL_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign PIO_LCD_CTRL_s1_any_bursting_master_saved_grant = 0;

  //PIO_LCD_CTRL_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign PIO_LCD_CTRL_s1_arb_share_counter_next_value = PIO_LCD_CTRL_s1_firsttransfer ? (PIO_LCD_CTRL_s1_arb_share_set_values - 1) : |PIO_LCD_CTRL_s1_arb_share_counter ? (PIO_LCD_CTRL_s1_arb_share_counter - 1) : 0;

  //PIO_LCD_CTRL_s1_allgrants all slave grants, which is an e_mux
  assign PIO_LCD_CTRL_s1_allgrants = |PIO_LCD_CTRL_s1_grant_vector;

  //PIO_LCD_CTRL_s1_end_xfer assignment, which is an e_assign
  assign PIO_LCD_CTRL_s1_end_xfer = ~(PIO_LCD_CTRL_s1_waits_for_read | PIO_LCD_CTRL_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_PIO_LCD_CTRL_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_PIO_LCD_CTRL_s1 = PIO_LCD_CTRL_s1_end_xfer & (~PIO_LCD_CTRL_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //PIO_LCD_CTRL_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign PIO_LCD_CTRL_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_PIO_LCD_CTRL_s1 & PIO_LCD_CTRL_s1_allgrants) | (end_xfer_arb_share_counter_term_PIO_LCD_CTRL_s1 & ~PIO_LCD_CTRL_s1_non_bursting_master_requests);

  //PIO_LCD_CTRL_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_CTRL_s1_arb_share_counter <= 0;
      else if (PIO_LCD_CTRL_s1_arb_counter_enable)
          PIO_LCD_CTRL_s1_arb_share_counter <= PIO_LCD_CTRL_s1_arb_share_counter_next_value;
    end


  //PIO_LCD_CTRL_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_CTRL_s1_slavearbiterlockenable <= 0;
      else if ((|PIO_LCD_CTRL_s1_master_qreq_vector & end_xfer_arb_share_counter_term_PIO_LCD_CTRL_s1) | (end_xfer_arb_share_counter_term_PIO_LCD_CTRL_s1 & ~PIO_LCD_CTRL_s1_non_bursting_master_requests))
          PIO_LCD_CTRL_s1_slavearbiterlockenable <= |PIO_LCD_CTRL_s1_arb_share_counter_next_value;
    end


  //cpu/data_master PIO_LCD_CTRL/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = PIO_LCD_CTRL_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //PIO_LCD_CTRL_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign PIO_LCD_CTRL_s1_slavearbiterlockenable2 = |PIO_LCD_CTRL_s1_arb_share_counter_next_value;

  //cpu/data_master PIO_LCD_CTRL/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = PIO_LCD_CTRL_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //PIO_LCD_CTRL_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign PIO_LCD_CTRL_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_PIO_LCD_CTRL_s1 = cpu_data_master_requests_PIO_LCD_CTRL_s1 & ~(((~cpu_data_master_waitrequest) & cpu_data_master_write));
  //PIO_LCD_CTRL_s1_writedata mux, which is an e_mux
  assign PIO_LCD_CTRL_s1_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_PIO_LCD_CTRL_s1 = cpu_data_master_qualified_request_PIO_LCD_CTRL_s1;

  //cpu/data_master saved-grant PIO_LCD_CTRL/s1, which is an e_assign
  assign cpu_data_master_saved_grant_PIO_LCD_CTRL_s1 = cpu_data_master_requests_PIO_LCD_CTRL_s1;

  //allow new arb cycle for PIO_LCD_CTRL/s1, which is an e_assign
  assign PIO_LCD_CTRL_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign PIO_LCD_CTRL_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign PIO_LCD_CTRL_s1_master_qreq_vector = 1;

  //PIO_LCD_CTRL_s1_reset_n assignment, which is an e_assign
  assign PIO_LCD_CTRL_s1_reset_n = reset_n;

  assign PIO_LCD_CTRL_s1_chipselect = cpu_data_master_granted_PIO_LCD_CTRL_s1;
  //PIO_LCD_CTRL_s1_firsttransfer first transaction, which is an e_assign
  assign PIO_LCD_CTRL_s1_firsttransfer = PIO_LCD_CTRL_s1_begins_xfer ? PIO_LCD_CTRL_s1_unreg_firsttransfer : PIO_LCD_CTRL_s1_reg_firsttransfer;

  //PIO_LCD_CTRL_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign PIO_LCD_CTRL_s1_unreg_firsttransfer = ~(PIO_LCD_CTRL_s1_slavearbiterlockenable & PIO_LCD_CTRL_s1_any_continuerequest);

  //PIO_LCD_CTRL_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_CTRL_s1_reg_firsttransfer <= 1'b1;
      else if (PIO_LCD_CTRL_s1_begins_xfer)
          PIO_LCD_CTRL_s1_reg_firsttransfer <= PIO_LCD_CTRL_s1_unreg_firsttransfer;
    end


  //PIO_LCD_CTRL_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign PIO_LCD_CTRL_s1_beginbursttransfer_internal = PIO_LCD_CTRL_s1_begins_xfer;

  //~PIO_LCD_CTRL_s1_write_n assignment, which is an e_mux
  assign PIO_LCD_CTRL_s1_write_n = ~(cpu_data_master_granted_PIO_LCD_CTRL_s1 & cpu_data_master_write);

  assign shifted_address_to_PIO_LCD_CTRL_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //PIO_LCD_CTRL_s1_address mux, which is an e_mux
  assign PIO_LCD_CTRL_s1_address = shifted_address_to_PIO_LCD_CTRL_s1_from_cpu_data_master >> 2;

  //d1_PIO_LCD_CTRL_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_PIO_LCD_CTRL_s1_end_xfer <= 1;
      else 
        d1_PIO_LCD_CTRL_s1_end_xfer <= PIO_LCD_CTRL_s1_end_xfer;
    end


  //PIO_LCD_CTRL_s1_waits_for_read in a cycle, which is an e_mux
  assign PIO_LCD_CTRL_s1_waits_for_read = PIO_LCD_CTRL_s1_in_a_read_cycle & PIO_LCD_CTRL_s1_begins_xfer;

  //PIO_LCD_CTRL_s1_in_a_read_cycle assignment, which is an e_assign
  assign PIO_LCD_CTRL_s1_in_a_read_cycle = cpu_data_master_granted_PIO_LCD_CTRL_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = PIO_LCD_CTRL_s1_in_a_read_cycle;

  //PIO_LCD_CTRL_s1_waits_for_write in a cycle, which is an e_mux
  assign PIO_LCD_CTRL_s1_waits_for_write = PIO_LCD_CTRL_s1_in_a_write_cycle & 0;

  //PIO_LCD_CTRL_s1_in_a_write_cycle assignment, which is an e_assign
  assign PIO_LCD_CTRL_s1_in_a_write_cycle = cpu_data_master_granted_PIO_LCD_CTRL_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = PIO_LCD_CTRL_s1_in_a_write_cycle;

  assign wait_for_PIO_LCD_CTRL_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //PIO_LCD_CTRL/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module PIO_LCD_G_s1_arbitrator (
                                 // inputs:
                                  PIO_LCD_G_s1_readdata,
                                  clk,
                                  cpu_data_master_address_to_slave,
                                  cpu_data_master_read,
                                  cpu_data_master_waitrequest,
                                  cpu_data_master_write,
                                  cpu_data_master_writedata,
                                  reset_n,

                                 // outputs:
                                  PIO_LCD_G_s1_address,
                                  PIO_LCD_G_s1_chipselect,
                                  PIO_LCD_G_s1_readdata_from_sa,
                                  PIO_LCD_G_s1_reset_n,
                                  PIO_LCD_G_s1_write_n,
                                  PIO_LCD_G_s1_writedata,
                                  cpu_data_master_granted_PIO_LCD_G_s1,
                                  cpu_data_master_qualified_request_PIO_LCD_G_s1,
                                  cpu_data_master_read_data_valid_PIO_LCD_G_s1,
                                  cpu_data_master_requests_PIO_LCD_G_s1,
                                  d1_PIO_LCD_G_s1_end_xfer
                               )
;

  output  [  1: 0] PIO_LCD_G_s1_address;
  output           PIO_LCD_G_s1_chipselect;
  output  [ 31: 0] PIO_LCD_G_s1_readdata_from_sa;
  output           PIO_LCD_G_s1_reset_n;
  output           PIO_LCD_G_s1_write_n;
  output  [ 31: 0] PIO_LCD_G_s1_writedata;
  output           cpu_data_master_granted_PIO_LCD_G_s1;
  output           cpu_data_master_qualified_request_PIO_LCD_G_s1;
  output           cpu_data_master_read_data_valid_PIO_LCD_G_s1;
  output           cpu_data_master_requests_PIO_LCD_G_s1;
  output           d1_PIO_LCD_G_s1_end_xfer;
  input   [ 31: 0] PIO_LCD_G_s1_readdata;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_read;
  input            cpu_data_master_waitrequest;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;

  wire    [  1: 0] PIO_LCD_G_s1_address;
  wire             PIO_LCD_G_s1_allgrants;
  wire             PIO_LCD_G_s1_allow_new_arb_cycle;
  wire             PIO_LCD_G_s1_any_bursting_master_saved_grant;
  wire             PIO_LCD_G_s1_any_continuerequest;
  wire             PIO_LCD_G_s1_arb_counter_enable;
  reg     [  1: 0] PIO_LCD_G_s1_arb_share_counter;
  wire    [  1: 0] PIO_LCD_G_s1_arb_share_counter_next_value;
  wire    [  1: 0] PIO_LCD_G_s1_arb_share_set_values;
  wire             PIO_LCD_G_s1_beginbursttransfer_internal;
  wire             PIO_LCD_G_s1_begins_xfer;
  wire             PIO_LCD_G_s1_chipselect;
  wire             PIO_LCD_G_s1_end_xfer;
  wire             PIO_LCD_G_s1_firsttransfer;
  wire             PIO_LCD_G_s1_grant_vector;
  wire             PIO_LCD_G_s1_in_a_read_cycle;
  wire             PIO_LCD_G_s1_in_a_write_cycle;
  wire             PIO_LCD_G_s1_master_qreq_vector;
  wire             PIO_LCD_G_s1_non_bursting_master_requests;
  wire    [ 31: 0] PIO_LCD_G_s1_readdata_from_sa;
  reg              PIO_LCD_G_s1_reg_firsttransfer;
  wire             PIO_LCD_G_s1_reset_n;
  reg              PIO_LCD_G_s1_slavearbiterlockenable;
  wire             PIO_LCD_G_s1_slavearbiterlockenable2;
  wire             PIO_LCD_G_s1_unreg_firsttransfer;
  wire             PIO_LCD_G_s1_waits_for_read;
  wire             PIO_LCD_G_s1_waits_for_write;
  wire             PIO_LCD_G_s1_write_n;
  wire    [ 31: 0] PIO_LCD_G_s1_writedata;
  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_PIO_LCD_G_s1;
  wire             cpu_data_master_qualified_request_PIO_LCD_G_s1;
  wire             cpu_data_master_read_data_valid_PIO_LCD_G_s1;
  wire             cpu_data_master_requests_PIO_LCD_G_s1;
  wire             cpu_data_master_saved_grant_PIO_LCD_G_s1;
  reg              d1_PIO_LCD_G_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_PIO_LCD_G_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 26: 0] shifted_address_to_PIO_LCD_G_s1_from_cpu_data_master;
  wire             wait_for_PIO_LCD_G_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~PIO_LCD_G_s1_end_xfer;
    end


  assign PIO_LCD_G_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_PIO_LCD_G_s1));
  //assign PIO_LCD_G_s1_readdata_from_sa = PIO_LCD_G_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign PIO_LCD_G_s1_readdata_from_sa = PIO_LCD_G_s1_readdata;

  assign cpu_data_master_requests_PIO_LCD_G_s1 = ({cpu_data_master_address_to_slave[26 : 4] , 4'b0} == 27'h1850) & (cpu_data_master_read | cpu_data_master_write);
  //PIO_LCD_G_s1_arb_share_counter set values, which is an e_mux
  assign PIO_LCD_G_s1_arb_share_set_values = 1;

  //PIO_LCD_G_s1_non_bursting_master_requests mux, which is an e_mux
  assign PIO_LCD_G_s1_non_bursting_master_requests = cpu_data_master_requests_PIO_LCD_G_s1;

  //PIO_LCD_G_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign PIO_LCD_G_s1_any_bursting_master_saved_grant = 0;

  //PIO_LCD_G_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign PIO_LCD_G_s1_arb_share_counter_next_value = PIO_LCD_G_s1_firsttransfer ? (PIO_LCD_G_s1_arb_share_set_values - 1) : |PIO_LCD_G_s1_arb_share_counter ? (PIO_LCD_G_s1_arb_share_counter - 1) : 0;

  //PIO_LCD_G_s1_allgrants all slave grants, which is an e_mux
  assign PIO_LCD_G_s1_allgrants = |PIO_LCD_G_s1_grant_vector;

  //PIO_LCD_G_s1_end_xfer assignment, which is an e_assign
  assign PIO_LCD_G_s1_end_xfer = ~(PIO_LCD_G_s1_waits_for_read | PIO_LCD_G_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_PIO_LCD_G_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_PIO_LCD_G_s1 = PIO_LCD_G_s1_end_xfer & (~PIO_LCD_G_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //PIO_LCD_G_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign PIO_LCD_G_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_PIO_LCD_G_s1 & PIO_LCD_G_s1_allgrants) | (end_xfer_arb_share_counter_term_PIO_LCD_G_s1 & ~PIO_LCD_G_s1_non_bursting_master_requests);

  //PIO_LCD_G_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_G_s1_arb_share_counter <= 0;
      else if (PIO_LCD_G_s1_arb_counter_enable)
          PIO_LCD_G_s1_arb_share_counter <= PIO_LCD_G_s1_arb_share_counter_next_value;
    end


  //PIO_LCD_G_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_G_s1_slavearbiterlockenable <= 0;
      else if ((|PIO_LCD_G_s1_master_qreq_vector & end_xfer_arb_share_counter_term_PIO_LCD_G_s1) | (end_xfer_arb_share_counter_term_PIO_LCD_G_s1 & ~PIO_LCD_G_s1_non_bursting_master_requests))
          PIO_LCD_G_s1_slavearbiterlockenable <= |PIO_LCD_G_s1_arb_share_counter_next_value;
    end


  //cpu/data_master PIO_LCD_G/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = PIO_LCD_G_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //PIO_LCD_G_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign PIO_LCD_G_s1_slavearbiterlockenable2 = |PIO_LCD_G_s1_arb_share_counter_next_value;

  //cpu/data_master PIO_LCD_G/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = PIO_LCD_G_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //PIO_LCD_G_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign PIO_LCD_G_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_PIO_LCD_G_s1 = cpu_data_master_requests_PIO_LCD_G_s1 & ~(((~cpu_data_master_waitrequest) & cpu_data_master_write));
  //PIO_LCD_G_s1_writedata mux, which is an e_mux
  assign PIO_LCD_G_s1_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_PIO_LCD_G_s1 = cpu_data_master_qualified_request_PIO_LCD_G_s1;

  //cpu/data_master saved-grant PIO_LCD_G/s1, which is an e_assign
  assign cpu_data_master_saved_grant_PIO_LCD_G_s1 = cpu_data_master_requests_PIO_LCD_G_s1;

  //allow new arb cycle for PIO_LCD_G/s1, which is an e_assign
  assign PIO_LCD_G_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign PIO_LCD_G_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign PIO_LCD_G_s1_master_qreq_vector = 1;

  //PIO_LCD_G_s1_reset_n assignment, which is an e_assign
  assign PIO_LCD_G_s1_reset_n = reset_n;

  assign PIO_LCD_G_s1_chipselect = cpu_data_master_granted_PIO_LCD_G_s1;
  //PIO_LCD_G_s1_firsttransfer first transaction, which is an e_assign
  assign PIO_LCD_G_s1_firsttransfer = PIO_LCD_G_s1_begins_xfer ? PIO_LCD_G_s1_unreg_firsttransfer : PIO_LCD_G_s1_reg_firsttransfer;

  //PIO_LCD_G_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign PIO_LCD_G_s1_unreg_firsttransfer = ~(PIO_LCD_G_s1_slavearbiterlockenable & PIO_LCD_G_s1_any_continuerequest);

  //PIO_LCD_G_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_G_s1_reg_firsttransfer <= 1'b1;
      else if (PIO_LCD_G_s1_begins_xfer)
          PIO_LCD_G_s1_reg_firsttransfer <= PIO_LCD_G_s1_unreg_firsttransfer;
    end


  //PIO_LCD_G_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign PIO_LCD_G_s1_beginbursttransfer_internal = PIO_LCD_G_s1_begins_xfer;

  //~PIO_LCD_G_s1_write_n assignment, which is an e_mux
  assign PIO_LCD_G_s1_write_n = ~(cpu_data_master_granted_PIO_LCD_G_s1 & cpu_data_master_write);

  assign shifted_address_to_PIO_LCD_G_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //PIO_LCD_G_s1_address mux, which is an e_mux
  assign PIO_LCD_G_s1_address = shifted_address_to_PIO_LCD_G_s1_from_cpu_data_master >> 2;

  //d1_PIO_LCD_G_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_PIO_LCD_G_s1_end_xfer <= 1;
      else 
        d1_PIO_LCD_G_s1_end_xfer <= PIO_LCD_G_s1_end_xfer;
    end


  //PIO_LCD_G_s1_waits_for_read in a cycle, which is an e_mux
  assign PIO_LCD_G_s1_waits_for_read = PIO_LCD_G_s1_in_a_read_cycle & PIO_LCD_G_s1_begins_xfer;

  //PIO_LCD_G_s1_in_a_read_cycle assignment, which is an e_assign
  assign PIO_LCD_G_s1_in_a_read_cycle = cpu_data_master_granted_PIO_LCD_G_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = PIO_LCD_G_s1_in_a_read_cycle;

  //PIO_LCD_G_s1_waits_for_write in a cycle, which is an e_mux
  assign PIO_LCD_G_s1_waits_for_write = PIO_LCD_G_s1_in_a_write_cycle & 0;

  //PIO_LCD_G_s1_in_a_write_cycle assignment, which is an e_assign
  assign PIO_LCD_G_s1_in_a_write_cycle = cpu_data_master_granted_PIO_LCD_G_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = PIO_LCD_G_s1_in_a_write_cycle;

  assign wait_for_PIO_LCD_G_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //PIO_LCD_G/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module PIO_LCD_PWM_s1_arbitrator (
                                   // inputs:
                                    PIO_LCD_PWM_s1_readdata,
                                    clk,
                                    cpu_data_master_address_to_slave,
                                    cpu_data_master_read,
                                    cpu_data_master_waitrequest,
                                    cpu_data_master_write,
                                    cpu_data_master_writedata,
                                    reset_n,

                                   // outputs:
                                    PIO_LCD_PWM_s1_address,
                                    PIO_LCD_PWM_s1_chipselect,
                                    PIO_LCD_PWM_s1_readdata_from_sa,
                                    PIO_LCD_PWM_s1_reset_n,
                                    PIO_LCD_PWM_s1_write_n,
                                    PIO_LCD_PWM_s1_writedata,
                                    cpu_data_master_granted_PIO_LCD_PWM_s1,
                                    cpu_data_master_qualified_request_PIO_LCD_PWM_s1,
                                    cpu_data_master_read_data_valid_PIO_LCD_PWM_s1,
                                    cpu_data_master_requests_PIO_LCD_PWM_s1,
                                    d1_PIO_LCD_PWM_s1_end_xfer
                                 )
;

  output  [  1: 0] PIO_LCD_PWM_s1_address;
  output           PIO_LCD_PWM_s1_chipselect;
  output  [ 31: 0] PIO_LCD_PWM_s1_readdata_from_sa;
  output           PIO_LCD_PWM_s1_reset_n;
  output           PIO_LCD_PWM_s1_write_n;
  output  [ 31: 0] PIO_LCD_PWM_s1_writedata;
  output           cpu_data_master_granted_PIO_LCD_PWM_s1;
  output           cpu_data_master_qualified_request_PIO_LCD_PWM_s1;
  output           cpu_data_master_read_data_valid_PIO_LCD_PWM_s1;
  output           cpu_data_master_requests_PIO_LCD_PWM_s1;
  output           d1_PIO_LCD_PWM_s1_end_xfer;
  input   [ 31: 0] PIO_LCD_PWM_s1_readdata;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_read;
  input            cpu_data_master_waitrequest;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;

  wire    [  1: 0] PIO_LCD_PWM_s1_address;
  wire             PIO_LCD_PWM_s1_allgrants;
  wire             PIO_LCD_PWM_s1_allow_new_arb_cycle;
  wire             PIO_LCD_PWM_s1_any_bursting_master_saved_grant;
  wire             PIO_LCD_PWM_s1_any_continuerequest;
  wire             PIO_LCD_PWM_s1_arb_counter_enable;
  reg     [  1: 0] PIO_LCD_PWM_s1_arb_share_counter;
  wire    [  1: 0] PIO_LCD_PWM_s1_arb_share_counter_next_value;
  wire    [  1: 0] PIO_LCD_PWM_s1_arb_share_set_values;
  wire             PIO_LCD_PWM_s1_beginbursttransfer_internal;
  wire             PIO_LCD_PWM_s1_begins_xfer;
  wire             PIO_LCD_PWM_s1_chipselect;
  wire             PIO_LCD_PWM_s1_end_xfer;
  wire             PIO_LCD_PWM_s1_firsttransfer;
  wire             PIO_LCD_PWM_s1_grant_vector;
  wire             PIO_LCD_PWM_s1_in_a_read_cycle;
  wire             PIO_LCD_PWM_s1_in_a_write_cycle;
  wire             PIO_LCD_PWM_s1_master_qreq_vector;
  wire             PIO_LCD_PWM_s1_non_bursting_master_requests;
  wire    [ 31: 0] PIO_LCD_PWM_s1_readdata_from_sa;
  reg              PIO_LCD_PWM_s1_reg_firsttransfer;
  wire             PIO_LCD_PWM_s1_reset_n;
  reg              PIO_LCD_PWM_s1_slavearbiterlockenable;
  wire             PIO_LCD_PWM_s1_slavearbiterlockenable2;
  wire             PIO_LCD_PWM_s1_unreg_firsttransfer;
  wire             PIO_LCD_PWM_s1_waits_for_read;
  wire             PIO_LCD_PWM_s1_waits_for_write;
  wire             PIO_LCD_PWM_s1_write_n;
  wire    [ 31: 0] PIO_LCD_PWM_s1_writedata;
  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_PIO_LCD_PWM_s1;
  wire             cpu_data_master_qualified_request_PIO_LCD_PWM_s1;
  wire             cpu_data_master_read_data_valid_PIO_LCD_PWM_s1;
  wire             cpu_data_master_requests_PIO_LCD_PWM_s1;
  wire             cpu_data_master_saved_grant_PIO_LCD_PWM_s1;
  reg              d1_PIO_LCD_PWM_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_PIO_LCD_PWM_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 26: 0] shifted_address_to_PIO_LCD_PWM_s1_from_cpu_data_master;
  wire             wait_for_PIO_LCD_PWM_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~PIO_LCD_PWM_s1_end_xfer;
    end


  assign PIO_LCD_PWM_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_PIO_LCD_PWM_s1));
  //assign PIO_LCD_PWM_s1_readdata_from_sa = PIO_LCD_PWM_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign PIO_LCD_PWM_s1_readdata_from_sa = PIO_LCD_PWM_s1_readdata;

  assign cpu_data_master_requests_PIO_LCD_PWM_s1 = ({cpu_data_master_address_to_slave[26 : 4] , 4'b0} == 27'h1820) & (cpu_data_master_read | cpu_data_master_write);
  //PIO_LCD_PWM_s1_arb_share_counter set values, which is an e_mux
  assign PIO_LCD_PWM_s1_arb_share_set_values = 1;

  //PIO_LCD_PWM_s1_non_bursting_master_requests mux, which is an e_mux
  assign PIO_LCD_PWM_s1_non_bursting_master_requests = cpu_data_master_requests_PIO_LCD_PWM_s1;

  //PIO_LCD_PWM_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign PIO_LCD_PWM_s1_any_bursting_master_saved_grant = 0;

  //PIO_LCD_PWM_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign PIO_LCD_PWM_s1_arb_share_counter_next_value = PIO_LCD_PWM_s1_firsttransfer ? (PIO_LCD_PWM_s1_arb_share_set_values - 1) : |PIO_LCD_PWM_s1_arb_share_counter ? (PIO_LCD_PWM_s1_arb_share_counter - 1) : 0;

  //PIO_LCD_PWM_s1_allgrants all slave grants, which is an e_mux
  assign PIO_LCD_PWM_s1_allgrants = |PIO_LCD_PWM_s1_grant_vector;

  //PIO_LCD_PWM_s1_end_xfer assignment, which is an e_assign
  assign PIO_LCD_PWM_s1_end_xfer = ~(PIO_LCD_PWM_s1_waits_for_read | PIO_LCD_PWM_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_PIO_LCD_PWM_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_PIO_LCD_PWM_s1 = PIO_LCD_PWM_s1_end_xfer & (~PIO_LCD_PWM_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //PIO_LCD_PWM_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign PIO_LCD_PWM_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_PIO_LCD_PWM_s1 & PIO_LCD_PWM_s1_allgrants) | (end_xfer_arb_share_counter_term_PIO_LCD_PWM_s1 & ~PIO_LCD_PWM_s1_non_bursting_master_requests);

  //PIO_LCD_PWM_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_PWM_s1_arb_share_counter <= 0;
      else if (PIO_LCD_PWM_s1_arb_counter_enable)
          PIO_LCD_PWM_s1_arb_share_counter <= PIO_LCD_PWM_s1_arb_share_counter_next_value;
    end


  //PIO_LCD_PWM_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_PWM_s1_slavearbiterlockenable <= 0;
      else if ((|PIO_LCD_PWM_s1_master_qreq_vector & end_xfer_arb_share_counter_term_PIO_LCD_PWM_s1) | (end_xfer_arb_share_counter_term_PIO_LCD_PWM_s1 & ~PIO_LCD_PWM_s1_non_bursting_master_requests))
          PIO_LCD_PWM_s1_slavearbiterlockenable <= |PIO_LCD_PWM_s1_arb_share_counter_next_value;
    end


  //cpu/data_master PIO_LCD_PWM/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = PIO_LCD_PWM_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //PIO_LCD_PWM_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign PIO_LCD_PWM_s1_slavearbiterlockenable2 = |PIO_LCD_PWM_s1_arb_share_counter_next_value;

  //cpu/data_master PIO_LCD_PWM/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = PIO_LCD_PWM_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //PIO_LCD_PWM_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign PIO_LCD_PWM_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_PIO_LCD_PWM_s1 = cpu_data_master_requests_PIO_LCD_PWM_s1 & ~(((~cpu_data_master_waitrequest) & cpu_data_master_write));
  //PIO_LCD_PWM_s1_writedata mux, which is an e_mux
  assign PIO_LCD_PWM_s1_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_PIO_LCD_PWM_s1 = cpu_data_master_qualified_request_PIO_LCD_PWM_s1;

  //cpu/data_master saved-grant PIO_LCD_PWM/s1, which is an e_assign
  assign cpu_data_master_saved_grant_PIO_LCD_PWM_s1 = cpu_data_master_requests_PIO_LCD_PWM_s1;

  //allow new arb cycle for PIO_LCD_PWM/s1, which is an e_assign
  assign PIO_LCD_PWM_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign PIO_LCD_PWM_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign PIO_LCD_PWM_s1_master_qreq_vector = 1;

  //PIO_LCD_PWM_s1_reset_n assignment, which is an e_assign
  assign PIO_LCD_PWM_s1_reset_n = reset_n;

  assign PIO_LCD_PWM_s1_chipselect = cpu_data_master_granted_PIO_LCD_PWM_s1;
  //PIO_LCD_PWM_s1_firsttransfer first transaction, which is an e_assign
  assign PIO_LCD_PWM_s1_firsttransfer = PIO_LCD_PWM_s1_begins_xfer ? PIO_LCD_PWM_s1_unreg_firsttransfer : PIO_LCD_PWM_s1_reg_firsttransfer;

  //PIO_LCD_PWM_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign PIO_LCD_PWM_s1_unreg_firsttransfer = ~(PIO_LCD_PWM_s1_slavearbiterlockenable & PIO_LCD_PWM_s1_any_continuerequest);

  //PIO_LCD_PWM_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_PWM_s1_reg_firsttransfer <= 1'b1;
      else if (PIO_LCD_PWM_s1_begins_xfer)
          PIO_LCD_PWM_s1_reg_firsttransfer <= PIO_LCD_PWM_s1_unreg_firsttransfer;
    end


  //PIO_LCD_PWM_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign PIO_LCD_PWM_s1_beginbursttransfer_internal = PIO_LCD_PWM_s1_begins_xfer;

  //~PIO_LCD_PWM_s1_write_n assignment, which is an e_mux
  assign PIO_LCD_PWM_s1_write_n = ~(cpu_data_master_granted_PIO_LCD_PWM_s1 & cpu_data_master_write);

  assign shifted_address_to_PIO_LCD_PWM_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //PIO_LCD_PWM_s1_address mux, which is an e_mux
  assign PIO_LCD_PWM_s1_address = shifted_address_to_PIO_LCD_PWM_s1_from_cpu_data_master >> 2;

  //d1_PIO_LCD_PWM_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_PIO_LCD_PWM_s1_end_xfer <= 1;
      else 
        d1_PIO_LCD_PWM_s1_end_xfer <= PIO_LCD_PWM_s1_end_xfer;
    end


  //PIO_LCD_PWM_s1_waits_for_read in a cycle, which is an e_mux
  assign PIO_LCD_PWM_s1_waits_for_read = PIO_LCD_PWM_s1_in_a_read_cycle & PIO_LCD_PWM_s1_begins_xfer;

  //PIO_LCD_PWM_s1_in_a_read_cycle assignment, which is an e_assign
  assign PIO_LCD_PWM_s1_in_a_read_cycle = cpu_data_master_granted_PIO_LCD_PWM_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = PIO_LCD_PWM_s1_in_a_read_cycle;

  //PIO_LCD_PWM_s1_waits_for_write in a cycle, which is an e_mux
  assign PIO_LCD_PWM_s1_waits_for_write = PIO_LCD_PWM_s1_in_a_write_cycle & 0;

  //PIO_LCD_PWM_s1_in_a_write_cycle assignment, which is an e_assign
  assign PIO_LCD_PWM_s1_in_a_write_cycle = cpu_data_master_granted_PIO_LCD_PWM_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = PIO_LCD_PWM_s1_in_a_write_cycle;

  assign wait_for_PIO_LCD_PWM_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //PIO_LCD_PWM/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module PIO_LCD_R_s1_arbitrator (
                                 // inputs:
                                  PIO_LCD_R_s1_readdata,
                                  clk,
                                  cpu_data_master_address_to_slave,
                                  cpu_data_master_read,
                                  cpu_data_master_waitrequest,
                                  cpu_data_master_write,
                                  cpu_data_master_writedata,
                                  reset_n,

                                 // outputs:
                                  PIO_LCD_R_s1_address,
                                  PIO_LCD_R_s1_chipselect,
                                  PIO_LCD_R_s1_readdata_from_sa,
                                  PIO_LCD_R_s1_reset_n,
                                  PIO_LCD_R_s1_write_n,
                                  PIO_LCD_R_s1_writedata,
                                  cpu_data_master_granted_PIO_LCD_R_s1,
                                  cpu_data_master_qualified_request_PIO_LCD_R_s1,
                                  cpu_data_master_read_data_valid_PIO_LCD_R_s1,
                                  cpu_data_master_requests_PIO_LCD_R_s1,
                                  d1_PIO_LCD_R_s1_end_xfer
                               )
;

  output  [  1: 0] PIO_LCD_R_s1_address;
  output           PIO_LCD_R_s1_chipselect;
  output  [ 31: 0] PIO_LCD_R_s1_readdata_from_sa;
  output           PIO_LCD_R_s1_reset_n;
  output           PIO_LCD_R_s1_write_n;
  output  [ 31: 0] PIO_LCD_R_s1_writedata;
  output           cpu_data_master_granted_PIO_LCD_R_s1;
  output           cpu_data_master_qualified_request_PIO_LCD_R_s1;
  output           cpu_data_master_read_data_valid_PIO_LCD_R_s1;
  output           cpu_data_master_requests_PIO_LCD_R_s1;
  output           d1_PIO_LCD_R_s1_end_xfer;
  input   [ 31: 0] PIO_LCD_R_s1_readdata;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_read;
  input            cpu_data_master_waitrequest;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;

  wire    [  1: 0] PIO_LCD_R_s1_address;
  wire             PIO_LCD_R_s1_allgrants;
  wire             PIO_LCD_R_s1_allow_new_arb_cycle;
  wire             PIO_LCD_R_s1_any_bursting_master_saved_grant;
  wire             PIO_LCD_R_s1_any_continuerequest;
  wire             PIO_LCD_R_s1_arb_counter_enable;
  reg     [  1: 0] PIO_LCD_R_s1_arb_share_counter;
  wire    [  1: 0] PIO_LCD_R_s1_arb_share_counter_next_value;
  wire    [  1: 0] PIO_LCD_R_s1_arb_share_set_values;
  wire             PIO_LCD_R_s1_beginbursttransfer_internal;
  wire             PIO_LCD_R_s1_begins_xfer;
  wire             PIO_LCD_R_s1_chipselect;
  wire             PIO_LCD_R_s1_end_xfer;
  wire             PIO_LCD_R_s1_firsttransfer;
  wire             PIO_LCD_R_s1_grant_vector;
  wire             PIO_LCD_R_s1_in_a_read_cycle;
  wire             PIO_LCD_R_s1_in_a_write_cycle;
  wire             PIO_LCD_R_s1_master_qreq_vector;
  wire             PIO_LCD_R_s1_non_bursting_master_requests;
  wire    [ 31: 0] PIO_LCD_R_s1_readdata_from_sa;
  reg              PIO_LCD_R_s1_reg_firsttransfer;
  wire             PIO_LCD_R_s1_reset_n;
  reg              PIO_LCD_R_s1_slavearbiterlockenable;
  wire             PIO_LCD_R_s1_slavearbiterlockenable2;
  wire             PIO_LCD_R_s1_unreg_firsttransfer;
  wire             PIO_LCD_R_s1_waits_for_read;
  wire             PIO_LCD_R_s1_waits_for_write;
  wire             PIO_LCD_R_s1_write_n;
  wire    [ 31: 0] PIO_LCD_R_s1_writedata;
  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_PIO_LCD_R_s1;
  wire             cpu_data_master_qualified_request_PIO_LCD_R_s1;
  wire             cpu_data_master_read_data_valid_PIO_LCD_R_s1;
  wire             cpu_data_master_requests_PIO_LCD_R_s1;
  wire             cpu_data_master_saved_grant_PIO_LCD_R_s1;
  reg              d1_PIO_LCD_R_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_PIO_LCD_R_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 26: 0] shifted_address_to_PIO_LCD_R_s1_from_cpu_data_master;
  wire             wait_for_PIO_LCD_R_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~PIO_LCD_R_s1_end_xfer;
    end


  assign PIO_LCD_R_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_PIO_LCD_R_s1));
  //assign PIO_LCD_R_s1_readdata_from_sa = PIO_LCD_R_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign PIO_LCD_R_s1_readdata_from_sa = PIO_LCD_R_s1_readdata;

  assign cpu_data_master_requests_PIO_LCD_R_s1 = ({cpu_data_master_address_to_slave[26 : 4] , 4'b0} == 27'h1860) & (cpu_data_master_read | cpu_data_master_write);
  //PIO_LCD_R_s1_arb_share_counter set values, which is an e_mux
  assign PIO_LCD_R_s1_arb_share_set_values = 1;

  //PIO_LCD_R_s1_non_bursting_master_requests mux, which is an e_mux
  assign PIO_LCD_R_s1_non_bursting_master_requests = cpu_data_master_requests_PIO_LCD_R_s1;

  //PIO_LCD_R_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign PIO_LCD_R_s1_any_bursting_master_saved_grant = 0;

  //PIO_LCD_R_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign PIO_LCD_R_s1_arb_share_counter_next_value = PIO_LCD_R_s1_firsttransfer ? (PIO_LCD_R_s1_arb_share_set_values - 1) : |PIO_LCD_R_s1_arb_share_counter ? (PIO_LCD_R_s1_arb_share_counter - 1) : 0;

  //PIO_LCD_R_s1_allgrants all slave grants, which is an e_mux
  assign PIO_LCD_R_s1_allgrants = |PIO_LCD_R_s1_grant_vector;

  //PIO_LCD_R_s1_end_xfer assignment, which is an e_assign
  assign PIO_LCD_R_s1_end_xfer = ~(PIO_LCD_R_s1_waits_for_read | PIO_LCD_R_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_PIO_LCD_R_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_PIO_LCD_R_s1 = PIO_LCD_R_s1_end_xfer & (~PIO_LCD_R_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //PIO_LCD_R_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign PIO_LCD_R_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_PIO_LCD_R_s1 & PIO_LCD_R_s1_allgrants) | (end_xfer_arb_share_counter_term_PIO_LCD_R_s1 & ~PIO_LCD_R_s1_non_bursting_master_requests);

  //PIO_LCD_R_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_R_s1_arb_share_counter <= 0;
      else if (PIO_LCD_R_s1_arb_counter_enable)
          PIO_LCD_R_s1_arb_share_counter <= PIO_LCD_R_s1_arb_share_counter_next_value;
    end


  //PIO_LCD_R_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_R_s1_slavearbiterlockenable <= 0;
      else if ((|PIO_LCD_R_s1_master_qreq_vector & end_xfer_arb_share_counter_term_PIO_LCD_R_s1) | (end_xfer_arb_share_counter_term_PIO_LCD_R_s1 & ~PIO_LCD_R_s1_non_bursting_master_requests))
          PIO_LCD_R_s1_slavearbiterlockenable <= |PIO_LCD_R_s1_arb_share_counter_next_value;
    end


  //cpu/data_master PIO_LCD_R/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = PIO_LCD_R_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //PIO_LCD_R_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign PIO_LCD_R_s1_slavearbiterlockenable2 = |PIO_LCD_R_s1_arb_share_counter_next_value;

  //cpu/data_master PIO_LCD_R/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = PIO_LCD_R_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //PIO_LCD_R_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign PIO_LCD_R_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_PIO_LCD_R_s1 = cpu_data_master_requests_PIO_LCD_R_s1 & ~(((~cpu_data_master_waitrequest) & cpu_data_master_write));
  //PIO_LCD_R_s1_writedata mux, which is an e_mux
  assign PIO_LCD_R_s1_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_PIO_LCD_R_s1 = cpu_data_master_qualified_request_PIO_LCD_R_s1;

  //cpu/data_master saved-grant PIO_LCD_R/s1, which is an e_assign
  assign cpu_data_master_saved_grant_PIO_LCD_R_s1 = cpu_data_master_requests_PIO_LCD_R_s1;

  //allow new arb cycle for PIO_LCD_R/s1, which is an e_assign
  assign PIO_LCD_R_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign PIO_LCD_R_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign PIO_LCD_R_s1_master_qreq_vector = 1;

  //PIO_LCD_R_s1_reset_n assignment, which is an e_assign
  assign PIO_LCD_R_s1_reset_n = reset_n;

  assign PIO_LCD_R_s1_chipselect = cpu_data_master_granted_PIO_LCD_R_s1;
  //PIO_LCD_R_s1_firsttransfer first transaction, which is an e_assign
  assign PIO_LCD_R_s1_firsttransfer = PIO_LCD_R_s1_begins_xfer ? PIO_LCD_R_s1_unreg_firsttransfer : PIO_LCD_R_s1_reg_firsttransfer;

  //PIO_LCD_R_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign PIO_LCD_R_s1_unreg_firsttransfer = ~(PIO_LCD_R_s1_slavearbiterlockenable & PIO_LCD_R_s1_any_continuerequest);

  //PIO_LCD_R_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LCD_R_s1_reg_firsttransfer <= 1'b1;
      else if (PIO_LCD_R_s1_begins_xfer)
          PIO_LCD_R_s1_reg_firsttransfer <= PIO_LCD_R_s1_unreg_firsttransfer;
    end


  //PIO_LCD_R_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign PIO_LCD_R_s1_beginbursttransfer_internal = PIO_LCD_R_s1_begins_xfer;

  //~PIO_LCD_R_s1_write_n assignment, which is an e_mux
  assign PIO_LCD_R_s1_write_n = ~(cpu_data_master_granted_PIO_LCD_R_s1 & cpu_data_master_write);

  assign shifted_address_to_PIO_LCD_R_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //PIO_LCD_R_s1_address mux, which is an e_mux
  assign PIO_LCD_R_s1_address = shifted_address_to_PIO_LCD_R_s1_from_cpu_data_master >> 2;

  //d1_PIO_LCD_R_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_PIO_LCD_R_s1_end_xfer <= 1;
      else 
        d1_PIO_LCD_R_s1_end_xfer <= PIO_LCD_R_s1_end_xfer;
    end


  //PIO_LCD_R_s1_waits_for_read in a cycle, which is an e_mux
  assign PIO_LCD_R_s1_waits_for_read = PIO_LCD_R_s1_in_a_read_cycle & PIO_LCD_R_s1_begins_xfer;

  //PIO_LCD_R_s1_in_a_read_cycle assignment, which is an e_assign
  assign PIO_LCD_R_s1_in_a_read_cycle = cpu_data_master_granted_PIO_LCD_R_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = PIO_LCD_R_s1_in_a_read_cycle;

  //PIO_LCD_R_s1_waits_for_write in a cycle, which is an e_mux
  assign PIO_LCD_R_s1_waits_for_write = PIO_LCD_R_s1_in_a_write_cycle & 0;

  //PIO_LCD_R_s1_in_a_write_cycle assignment, which is an e_assign
  assign PIO_LCD_R_s1_in_a_write_cycle = cpu_data_master_granted_PIO_LCD_R_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = PIO_LCD_R_s1_in_a_write_cycle;

  assign wait_for_PIO_LCD_R_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //PIO_LCD_R/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module PIO_LED_s1_arbitrator (
                               // inputs:
                                PIO_LED_s1_readdata,
                                clk,
                                cpu_data_master_address_to_slave,
                                cpu_data_master_read,
                                cpu_data_master_waitrequest,
                                cpu_data_master_write,
                                cpu_data_master_writedata,
                                reset_n,

                               // outputs:
                                PIO_LED_s1_address,
                                PIO_LED_s1_chipselect,
                                PIO_LED_s1_readdata_from_sa,
                                PIO_LED_s1_reset_n,
                                PIO_LED_s1_write_n,
                                PIO_LED_s1_writedata,
                                cpu_data_master_granted_PIO_LED_s1,
                                cpu_data_master_qualified_request_PIO_LED_s1,
                                cpu_data_master_read_data_valid_PIO_LED_s1,
                                cpu_data_master_requests_PIO_LED_s1,
                                d1_PIO_LED_s1_end_xfer
                             )
;

  output  [  1: 0] PIO_LED_s1_address;
  output           PIO_LED_s1_chipselect;
  output  [ 31: 0] PIO_LED_s1_readdata_from_sa;
  output           PIO_LED_s1_reset_n;
  output           PIO_LED_s1_write_n;
  output  [ 31: 0] PIO_LED_s1_writedata;
  output           cpu_data_master_granted_PIO_LED_s1;
  output           cpu_data_master_qualified_request_PIO_LED_s1;
  output           cpu_data_master_read_data_valid_PIO_LED_s1;
  output           cpu_data_master_requests_PIO_LED_s1;
  output           d1_PIO_LED_s1_end_xfer;
  input   [ 31: 0] PIO_LED_s1_readdata;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_read;
  input            cpu_data_master_waitrequest;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;

  wire    [  1: 0] PIO_LED_s1_address;
  wire             PIO_LED_s1_allgrants;
  wire             PIO_LED_s1_allow_new_arb_cycle;
  wire             PIO_LED_s1_any_bursting_master_saved_grant;
  wire             PIO_LED_s1_any_continuerequest;
  wire             PIO_LED_s1_arb_counter_enable;
  reg     [  1: 0] PIO_LED_s1_arb_share_counter;
  wire    [  1: 0] PIO_LED_s1_arb_share_counter_next_value;
  wire    [  1: 0] PIO_LED_s1_arb_share_set_values;
  wire             PIO_LED_s1_beginbursttransfer_internal;
  wire             PIO_LED_s1_begins_xfer;
  wire             PIO_LED_s1_chipselect;
  wire             PIO_LED_s1_end_xfer;
  wire             PIO_LED_s1_firsttransfer;
  wire             PIO_LED_s1_grant_vector;
  wire             PIO_LED_s1_in_a_read_cycle;
  wire             PIO_LED_s1_in_a_write_cycle;
  wire             PIO_LED_s1_master_qreq_vector;
  wire             PIO_LED_s1_non_bursting_master_requests;
  wire    [ 31: 0] PIO_LED_s1_readdata_from_sa;
  reg              PIO_LED_s1_reg_firsttransfer;
  wire             PIO_LED_s1_reset_n;
  reg              PIO_LED_s1_slavearbiterlockenable;
  wire             PIO_LED_s1_slavearbiterlockenable2;
  wire             PIO_LED_s1_unreg_firsttransfer;
  wire             PIO_LED_s1_waits_for_read;
  wire             PIO_LED_s1_waits_for_write;
  wire             PIO_LED_s1_write_n;
  wire    [ 31: 0] PIO_LED_s1_writedata;
  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_PIO_LED_s1;
  wire             cpu_data_master_qualified_request_PIO_LED_s1;
  wire             cpu_data_master_read_data_valid_PIO_LED_s1;
  wire             cpu_data_master_requests_PIO_LED_s1;
  wire             cpu_data_master_saved_grant_PIO_LED_s1;
  reg              d1_PIO_LED_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_PIO_LED_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 26: 0] shifted_address_to_PIO_LED_s1_from_cpu_data_master;
  wire             wait_for_PIO_LED_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~PIO_LED_s1_end_xfer;
    end


  assign PIO_LED_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_PIO_LED_s1));
  //assign PIO_LED_s1_readdata_from_sa = PIO_LED_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign PIO_LED_s1_readdata_from_sa = PIO_LED_s1_readdata;

  assign cpu_data_master_requests_PIO_LED_s1 = ({cpu_data_master_address_to_slave[26 : 4] , 4'b0} == 27'h1880) & (cpu_data_master_read | cpu_data_master_write);
  //PIO_LED_s1_arb_share_counter set values, which is an e_mux
  assign PIO_LED_s1_arb_share_set_values = 1;

  //PIO_LED_s1_non_bursting_master_requests mux, which is an e_mux
  assign PIO_LED_s1_non_bursting_master_requests = cpu_data_master_requests_PIO_LED_s1;

  //PIO_LED_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign PIO_LED_s1_any_bursting_master_saved_grant = 0;

  //PIO_LED_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign PIO_LED_s1_arb_share_counter_next_value = PIO_LED_s1_firsttransfer ? (PIO_LED_s1_arb_share_set_values - 1) : |PIO_LED_s1_arb_share_counter ? (PIO_LED_s1_arb_share_counter - 1) : 0;

  //PIO_LED_s1_allgrants all slave grants, which is an e_mux
  assign PIO_LED_s1_allgrants = |PIO_LED_s1_grant_vector;

  //PIO_LED_s1_end_xfer assignment, which is an e_assign
  assign PIO_LED_s1_end_xfer = ~(PIO_LED_s1_waits_for_read | PIO_LED_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_PIO_LED_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_PIO_LED_s1 = PIO_LED_s1_end_xfer & (~PIO_LED_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //PIO_LED_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign PIO_LED_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_PIO_LED_s1 & PIO_LED_s1_allgrants) | (end_xfer_arb_share_counter_term_PIO_LED_s1 & ~PIO_LED_s1_non_bursting_master_requests);

  //PIO_LED_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LED_s1_arb_share_counter <= 0;
      else if (PIO_LED_s1_arb_counter_enable)
          PIO_LED_s1_arb_share_counter <= PIO_LED_s1_arb_share_counter_next_value;
    end


  //PIO_LED_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LED_s1_slavearbiterlockenable <= 0;
      else if ((|PIO_LED_s1_master_qreq_vector & end_xfer_arb_share_counter_term_PIO_LED_s1) | (end_xfer_arb_share_counter_term_PIO_LED_s1 & ~PIO_LED_s1_non_bursting_master_requests))
          PIO_LED_s1_slavearbiterlockenable <= |PIO_LED_s1_arb_share_counter_next_value;
    end


  //cpu/data_master PIO_LED/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = PIO_LED_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //PIO_LED_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign PIO_LED_s1_slavearbiterlockenable2 = |PIO_LED_s1_arb_share_counter_next_value;

  //cpu/data_master PIO_LED/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = PIO_LED_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //PIO_LED_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign PIO_LED_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_PIO_LED_s1 = cpu_data_master_requests_PIO_LED_s1 & ~(((~cpu_data_master_waitrequest) & cpu_data_master_write));
  //PIO_LED_s1_writedata mux, which is an e_mux
  assign PIO_LED_s1_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_PIO_LED_s1 = cpu_data_master_qualified_request_PIO_LED_s1;

  //cpu/data_master saved-grant PIO_LED/s1, which is an e_assign
  assign cpu_data_master_saved_grant_PIO_LED_s1 = cpu_data_master_requests_PIO_LED_s1;

  //allow new arb cycle for PIO_LED/s1, which is an e_assign
  assign PIO_LED_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign PIO_LED_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign PIO_LED_s1_master_qreq_vector = 1;

  //PIO_LED_s1_reset_n assignment, which is an e_assign
  assign PIO_LED_s1_reset_n = reset_n;

  assign PIO_LED_s1_chipselect = cpu_data_master_granted_PIO_LED_s1;
  //PIO_LED_s1_firsttransfer first transaction, which is an e_assign
  assign PIO_LED_s1_firsttransfer = PIO_LED_s1_begins_xfer ? PIO_LED_s1_unreg_firsttransfer : PIO_LED_s1_reg_firsttransfer;

  //PIO_LED_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign PIO_LED_s1_unreg_firsttransfer = ~(PIO_LED_s1_slavearbiterlockenable & PIO_LED_s1_any_continuerequest);

  //PIO_LED_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          PIO_LED_s1_reg_firsttransfer <= 1'b1;
      else if (PIO_LED_s1_begins_xfer)
          PIO_LED_s1_reg_firsttransfer <= PIO_LED_s1_unreg_firsttransfer;
    end


  //PIO_LED_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign PIO_LED_s1_beginbursttransfer_internal = PIO_LED_s1_begins_xfer;

  //~PIO_LED_s1_write_n assignment, which is an e_mux
  assign PIO_LED_s1_write_n = ~(cpu_data_master_granted_PIO_LED_s1 & cpu_data_master_write);

  assign shifted_address_to_PIO_LED_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //PIO_LED_s1_address mux, which is an e_mux
  assign PIO_LED_s1_address = shifted_address_to_PIO_LED_s1_from_cpu_data_master >> 2;

  //d1_PIO_LED_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_PIO_LED_s1_end_xfer <= 1;
      else 
        d1_PIO_LED_s1_end_xfer <= PIO_LED_s1_end_xfer;
    end


  //PIO_LED_s1_waits_for_read in a cycle, which is an e_mux
  assign PIO_LED_s1_waits_for_read = PIO_LED_s1_in_a_read_cycle & PIO_LED_s1_begins_xfer;

  //PIO_LED_s1_in_a_read_cycle assignment, which is an e_assign
  assign PIO_LED_s1_in_a_read_cycle = cpu_data_master_granted_PIO_LED_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = PIO_LED_s1_in_a_read_cycle;

  //PIO_LED_s1_waits_for_write in a cycle, which is an e_mux
  assign PIO_LED_s1_waits_for_write = PIO_LED_s1_in_a_write_cycle & 0;

  //PIO_LED_s1_in_a_write_cycle assignment, which is an e_assign
  assign PIO_LED_s1_in_a_write_cycle = cpu_data_master_granted_PIO_LED_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = PIO_LED_s1_in_a_write_cycle;

  assign wait_for_PIO_LED_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //PIO_LED/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module RS232_s1_arbitrator (
                             // inputs:
                              RS232_s1_dataavailable,
                              RS232_s1_irq,
                              RS232_s1_readdata,
                              RS232_s1_readyfordata,
                              clk,
                              cpu_data_master_address_to_slave,
                              cpu_data_master_read,
                              cpu_data_master_write,
                              cpu_data_master_writedata,
                              reset_n,

                             // outputs:
                              RS232_s1_address,
                              RS232_s1_begintransfer,
                              RS232_s1_chipselect,
                              RS232_s1_dataavailable_from_sa,
                              RS232_s1_irq_from_sa,
                              RS232_s1_read_n,
                              RS232_s1_readdata_from_sa,
                              RS232_s1_readyfordata_from_sa,
                              RS232_s1_reset_n,
                              RS232_s1_write_n,
                              RS232_s1_writedata,
                              cpu_data_master_granted_RS232_s1,
                              cpu_data_master_qualified_request_RS232_s1,
                              cpu_data_master_read_data_valid_RS232_s1,
                              cpu_data_master_requests_RS232_s1,
                              d1_RS232_s1_end_xfer
                           )
;

  output  [  2: 0] RS232_s1_address;
  output           RS232_s1_begintransfer;
  output           RS232_s1_chipselect;
  output           RS232_s1_dataavailable_from_sa;
  output           RS232_s1_irq_from_sa;
  output           RS232_s1_read_n;
  output  [ 15: 0] RS232_s1_readdata_from_sa;
  output           RS232_s1_readyfordata_from_sa;
  output           RS232_s1_reset_n;
  output           RS232_s1_write_n;
  output  [ 15: 0] RS232_s1_writedata;
  output           cpu_data_master_granted_RS232_s1;
  output           cpu_data_master_qualified_request_RS232_s1;
  output           cpu_data_master_read_data_valid_RS232_s1;
  output           cpu_data_master_requests_RS232_s1;
  output           d1_RS232_s1_end_xfer;
  input            RS232_s1_dataavailable;
  input            RS232_s1_irq;
  input   [ 15: 0] RS232_s1_readdata;
  input            RS232_s1_readyfordata;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_read;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;

  wire    [  2: 0] RS232_s1_address;
  wire             RS232_s1_allgrants;
  wire             RS232_s1_allow_new_arb_cycle;
  wire             RS232_s1_any_bursting_master_saved_grant;
  wire             RS232_s1_any_continuerequest;
  wire             RS232_s1_arb_counter_enable;
  reg     [  1: 0] RS232_s1_arb_share_counter;
  wire    [  1: 0] RS232_s1_arb_share_counter_next_value;
  wire    [  1: 0] RS232_s1_arb_share_set_values;
  wire             RS232_s1_beginbursttransfer_internal;
  wire             RS232_s1_begins_xfer;
  wire             RS232_s1_begintransfer;
  wire             RS232_s1_chipselect;
  wire             RS232_s1_dataavailable_from_sa;
  wire             RS232_s1_end_xfer;
  wire             RS232_s1_firsttransfer;
  wire             RS232_s1_grant_vector;
  wire             RS232_s1_in_a_read_cycle;
  wire             RS232_s1_in_a_write_cycle;
  wire             RS232_s1_irq_from_sa;
  wire             RS232_s1_master_qreq_vector;
  wire             RS232_s1_non_bursting_master_requests;
  wire             RS232_s1_read_n;
  wire    [ 15: 0] RS232_s1_readdata_from_sa;
  wire             RS232_s1_readyfordata_from_sa;
  reg              RS232_s1_reg_firsttransfer;
  wire             RS232_s1_reset_n;
  reg              RS232_s1_slavearbiterlockenable;
  wire             RS232_s1_slavearbiterlockenable2;
  wire             RS232_s1_unreg_firsttransfer;
  wire             RS232_s1_waits_for_read;
  wire             RS232_s1_waits_for_write;
  wire             RS232_s1_write_n;
  wire    [ 15: 0] RS232_s1_writedata;
  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_RS232_s1;
  wire             cpu_data_master_qualified_request_RS232_s1;
  wire             cpu_data_master_read_data_valid_RS232_s1;
  wire             cpu_data_master_requests_RS232_s1;
  wire             cpu_data_master_saved_grant_RS232_s1;
  reg              d1_RS232_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_RS232_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 26: 0] shifted_address_to_RS232_s1_from_cpu_data_master;
  wire             wait_for_RS232_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~RS232_s1_end_xfer;
    end


  assign RS232_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_RS232_s1));
  //assign RS232_s1_readdata_from_sa = RS232_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign RS232_s1_readdata_from_sa = RS232_s1_readdata;

  assign cpu_data_master_requests_RS232_s1 = ({cpu_data_master_address_to_slave[26 : 5] , 5'b0} == 27'h1800) & (cpu_data_master_read | cpu_data_master_write);
  //assign RS232_s1_dataavailable_from_sa = RS232_s1_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign RS232_s1_dataavailable_from_sa = RS232_s1_dataavailable;

  //assign RS232_s1_readyfordata_from_sa = RS232_s1_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign RS232_s1_readyfordata_from_sa = RS232_s1_readyfordata;

  //RS232_s1_arb_share_counter set values, which is an e_mux
  assign RS232_s1_arb_share_set_values = 1;

  //RS232_s1_non_bursting_master_requests mux, which is an e_mux
  assign RS232_s1_non_bursting_master_requests = cpu_data_master_requests_RS232_s1;

  //RS232_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign RS232_s1_any_bursting_master_saved_grant = 0;

  //RS232_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign RS232_s1_arb_share_counter_next_value = RS232_s1_firsttransfer ? (RS232_s1_arb_share_set_values - 1) : |RS232_s1_arb_share_counter ? (RS232_s1_arb_share_counter - 1) : 0;

  //RS232_s1_allgrants all slave grants, which is an e_mux
  assign RS232_s1_allgrants = |RS232_s1_grant_vector;

  //RS232_s1_end_xfer assignment, which is an e_assign
  assign RS232_s1_end_xfer = ~(RS232_s1_waits_for_read | RS232_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_RS232_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_RS232_s1 = RS232_s1_end_xfer & (~RS232_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //RS232_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign RS232_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_RS232_s1 & RS232_s1_allgrants) | (end_xfer_arb_share_counter_term_RS232_s1 & ~RS232_s1_non_bursting_master_requests);

  //RS232_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          RS232_s1_arb_share_counter <= 0;
      else if (RS232_s1_arb_counter_enable)
          RS232_s1_arb_share_counter <= RS232_s1_arb_share_counter_next_value;
    end


  //RS232_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          RS232_s1_slavearbiterlockenable <= 0;
      else if ((|RS232_s1_master_qreq_vector & end_xfer_arb_share_counter_term_RS232_s1) | (end_xfer_arb_share_counter_term_RS232_s1 & ~RS232_s1_non_bursting_master_requests))
          RS232_s1_slavearbiterlockenable <= |RS232_s1_arb_share_counter_next_value;
    end


  //cpu/data_master RS232/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = RS232_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //RS232_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign RS232_s1_slavearbiterlockenable2 = |RS232_s1_arb_share_counter_next_value;

  //cpu/data_master RS232/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = RS232_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //RS232_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign RS232_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_RS232_s1 = cpu_data_master_requests_RS232_s1;
  //RS232_s1_writedata mux, which is an e_mux
  assign RS232_s1_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_RS232_s1 = cpu_data_master_qualified_request_RS232_s1;

  //cpu/data_master saved-grant RS232/s1, which is an e_assign
  assign cpu_data_master_saved_grant_RS232_s1 = cpu_data_master_requests_RS232_s1;

  //allow new arb cycle for RS232/s1, which is an e_assign
  assign RS232_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign RS232_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign RS232_s1_master_qreq_vector = 1;

  assign RS232_s1_begintransfer = RS232_s1_begins_xfer;
  //RS232_s1_reset_n assignment, which is an e_assign
  assign RS232_s1_reset_n = reset_n;

  assign RS232_s1_chipselect = cpu_data_master_granted_RS232_s1;
  //RS232_s1_firsttransfer first transaction, which is an e_assign
  assign RS232_s1_firsttransfer = RS232_s1_begins_xfer ? RS232_s1_unreg_firsttransfer : RS232_s1_reg_firsttransfer;

  //RS232_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign RS232_s1_unreg_firsttransfer = ~(RS232_s1_slavearbiterlockenable & RS232_s1_any_continuerequest);

  //RS232_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          RS232_s1_reg_firsttransfer <= 1'b1;
      else if (RS232_s1_begins_xfer)
          RS232_s1_reg_firsttransfer <= RS232_s1_unreg_firsttransfer;
    end


  //RS232_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign RS232_s1_beginbursttransfer_internal = RS232_s1_begins_xfer;

  //~RS232_s1_read_n assignment, which is an e_mux
  assign RS232_s1_read_n = ~(cpu_data_master_granted_RS232_s1 & cpu_data_master_read);

  //~RS232_s1_write_n assignment, which is an e_mux
  assign RS232_s1_write_n = ~(cpu_data_master_granted_RS232_s1 & cpu_data_master_write);

  assign shifted_address_to_RS232_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //RS232_s1_address mux, which is an e_mux
  assign RS232_s1_address = shifted_address_to_RS232_s1_from_cpu_data_master >> 2;

  //d1_RS232_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_RS232_s1_end_xfer <= 1;
      else 
        d1_RS232_s1_end_xfer <= RS232_s1_end_xfer;
    end


  //RS232_s1_waits_for_read in a cycle, which is an e_mux
  assign RS232_s1_waits_for_read = RS232_s1_in_a_read_cycle & RS232_s1_begins_xfer;

  //RS232_s1_in_a_read_cycle assignment, which is an e_assign
  assign RS232_s1_in_a_read_cycle = cpu_data_master_granted_RS232_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = RS232_s1_in_a_read_cycle;

  //RS232_s1_waits_for_write in a cycle, which is an e_mux
  assign RS232_s1_waits_for_write = RS232_s1_in_a_write_cycle & RS232_s1_begins_xfer;

  //RS232_s1_in_a_write_cycle assignment, which is an e_assign
  assign RS232_s1_in_a_write_cycle = cpu_data_master_granted_RS232_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = RS232_s1_in_a_write_cycle;

  assign wait_for_RS232_s1_counter = 0;
  //assign RS232_s1_irq_from_sa = RS232_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign RS232_s1_irq_from_sa = RS232_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //RS232/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_jtag_debug_module_arbitrator (
                                          // inputs:
                                           clk,
                                           cpu_data_master_address_to_slave,
                                           cpu_data_master_byteenable,
                                           cpu_data_master_debugaccess,
                                           cpu_data_master_read,
                                           cpu_data_master_waitrequest,
                                           cpu_data_master_write,
                                           cpu_data_master_writedata,
                                           cpu_instruction_master_address_to_slave,
                                           cpu_instruction_master_latency_counter,
                                           cpu_instruction_master_read,
                                           cpu_instruction_master_read_data_valid_sdram_s1_shift_register,
                                           cpu_jtag_debug_module_readdata,
                                           cpu_jtag_debug_module_resetrequest,
                                           reset_n,

                                          // outputs:
                                           cpu_data_master_granted_cpu_jtag_debug_module,
                                           cpu_data_master_qualified_request_cpu_jtag_debug_module,
                                           cpu_data_master_read_data_valid_cpu_jtag_debug_module,
                                           cpu_data_master_requests_cpu_jtag_debug_module,
                                           cpu_instruction_master_granted_cpu_jtag_debug_module,
                                           cpu_instruction_master_qualified_request_cpu_jtag_debug_module,
                                           cpu_instruction_master_read_data_valid_cpu_jtag_debug_module,
                                           cpu_instruction_master_requests_cpu_jtag_debug_module,
                                           cpu_jtag_debug_module_address,
                                           cpu_jtag_debug_module_begintransfer,
                                           cpu_jtag_debug_module_byteenable,
                                           cpu_jtag_debug_module_chipselect,
                                           cpu_jtag_debug_module_debugaccess,
                                           cpu_jtag_debug_module_readdata_from_sa,
                                           cpu_jtag_debug_module_reset_n,
                                           cpu_jtag_debug_module_resetrequest_from_sa,
                                           cpu_jtag_debug_module_write,
                                           cpu_jtag_debug_module_writedata,
                                           d1_cpu_jtag_debug_module_end_xfer
                                        )
;

  output           cpu_data_master_granted_cpu_jtag_debug_module;
  output           cpu_data_master_qualified_request_cpu_jtag_debug_module;
  output           cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  output           cpu_data_master_requests_cpu_jtag_debug_module;
  output           cpu_instruction_master_granted_cpu_jtag_debug_module;
  output           cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  output           cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  output           cpu_instruction_master_requests_cpu_jtag_debug_module;
  output  [  8: 0] cpu_jtag_debug_module_address;
  output           cpu_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_jtag_debug_module_byteenable;
  output           cpu_jtag_debug_module_chipselect;
  output           cpu_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  output           cpu_jtag_debug_module_reset_n;
  output           cpu_jtag_debug_module_resetrequest_from_sa;
  output           cpu_jtag_debug_module_write;
  output  [ 31: 0] cpu_jtag_debug_module_writedata;
  output           d1_cpu_jtag_debug_module_end_xfer;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_read;
  input            cpu_data_master_waitrequest;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 26: 0] cpu_instruction_master_address_to_slave;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_sdram_s1_shift_register;
  input   [ 31: 0] cpu_jtag_debug_module_readdata;
  input            cpu_jtag_debug_module_resetrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_cpu_jtag_debug_module;
  wire             cpu_data_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_data_master_requests_cpu_jtag_debug_module;
  wire             cpu_data_master_saved_grant_cpu_jtag_debug_module;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_cpu_jtag_debug_module;
  wire             cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_instruction_master_requests_cpu_jtag_debug_module;
  wire             cpu_instruction_master_saved_grant_cpu_jtag_debug_module;
  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_allgrants;
  wire             cpu_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_jtag_debug_module_any_continuerequest;
  reg     [  1: 0] cpu_jtag_debug_module_arb_addend;
  wire             cpu_jtag_debug_module_arb_counter_enable;
  reg     [  1: 0] cpu_jtag_debug_module_arb_share_counter;
  wire    [  1: 0] cpu_jtag_debug_module_arb_share_counter_next_value;
  wire    [  1: 0] cpu_jtag_debug_module_arb_share_set_values;
  wire    [  1: 0] cpu_jtag_debug_module_arb_winner;
  wire             cpu_jtag_debug_module_arbitration_holdoff_internal;
  wire             cpu_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_jtag_debug_module_begins_xfer;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire    [  3: 0] cpu_jtag_debug_module_chosen_master_double_vector;
  wire    [  1: 0] cpu_jtag_debug_module_chosen_master_rot_left;
  wire             cpu_jtag_debug_module_debugaccess;
  wire             cpu_jtag_debug_module_end_xfer;
  wire             cpu_jtag_debug_module_firsttransfer;
  wire    [  1: 0] cpu_jtag_debug_module_grant_vector;
  wire             cpu_jtag_debug_module_in_a_read_cycle;
  wire             cpu_jtag_debug_module_in_a_write_cycle;
  wire    [  1: 0] cpu_jtag_debug_module_master_qreq_vector;
  wire             cpu_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  reg              cpu_jtag_debug_module_reg_firsttransfer;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  reg     [  1: 0] cpu_jtag_debug_module_saved_chosen_master_vector;
  reg              cpu_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_jtag_debug_module_waits_for_read;
  wire             cpu_jtag_debug_module_waits_for_write;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  reg              d1_cpu_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module;
  reg              last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module;
  wire    [ 26: 0] shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master;
  wire    [ 26: 0] shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master;
  wire             wait_for_cpu_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_jtag_debug_module_end_xfer;
    end


  assign cpu_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_cpu_jtag_debug_module | cpu_instruction_master_qualified_request_cpu_jtag_debug_module));
  //assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata;

  assign cpu_data_master_requests_cpu_jtag_debug_module = ({cpu_data_master_address_to_slave[26 : 11] , 11'b0} == 27'h1000) & (cpu_data_master_read | cpu_data_master_write);
  //cpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_jtag_debug_module_arb_share_set_values = 1;

  //cpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_jtag_debug_module_non_bursting_master_requests = cpu_data_master_requests_cpu_jtag_debug_module |
    cpu_instruction_master_requests_cpu_jtag_debug_module |
    cpu_data_master_requests_cpu_jtag_debug_module |
    cpu_instruction_master_requests_cpu_jtag_debug_module;

  //cpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_jtag_debug_module_any_bursting_master_saved_grant = 0;

  //cpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_jtag_debug_module_arb_share_counter_next_value = cpu_jtag_debug_module_firsttransfer ? (cpu_jtag_debug_module_arb_share_set_values - 1) : |cpu_jtag_debug_module_arb_share_counter ? (cpu_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_jtag_debug_module_allgrants = (|cpu_jtag_debug_module_grant_vector) |
    (|cpu_jtag_debug_module_grant_vector) |
    (|cpu_jtag_debug_module_grant_vector) |
    (|cpu_jtag_debug_module_grant_vector);

  //cpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_jtag_debug_module_end_xfer = ~(cpu_jtag_debug_module_waits_for_read | cpu_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_jtag_debug_module = cpu_jtag_debug_module_end_xfer & (~cpu_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & cpu_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests);

  //cpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_jtag_debug_module_arb_counter_enable)
          cpu_jtag_debug_module_arb_share_counter <= cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests))
          cpu_jtag_debug_module_slavearbiterlockenable <= |cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu/data_master cpu/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = cpu_jtag_debug_module_slavearbiterlockenable & cpu_data_master_continuerequest;

  //cpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_jtag_debug_module_slavearbiterlockenable2 = |cpu_jtag_debug_module_arb_share_counter_next_value;

  //cpu/data_master cpu/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = cpu_jtag_debug_module_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master cpu/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = cpu_jtag_debug_module_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master cpu/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = cpu_jtag_debug_module_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted cpu/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module <= cpu_instruction_master_saved_grant_cpu_jtag_debug_module ? 1 : (cpu_jtag_debug_module_arbitration_holdoff_internal | ~cpu_instruction_master_requests_cpu_jtag_debug_module) ? 0 : last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module & cpu_instruction_master_requests_cpu_jtag_debug_module;

  //cpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  assign cpu_jtag_debug_module_any_continuerequest = cpu_instruction_master_continuerequest |
    cpu_data_master_continuerequest;

  assign cpu_data_master_qualified_request_cpu_jtag_debug_module = cpu_data_master_requests_cpu_jtag_debug_module & ~(((~cpu_data_master_waitrequest) & cpu_data_master_write) | cpu_instruction_master_arbiterlock);
  //cpu_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_jtag_debug_module_writedata = cpu_data_master_writedata;

  assign cpu_instruction_master_requests_cpu_jtag_debug_module = (({cpu_instruction_master_address_to_slave[26 : 11] , 11'b0} == 27'h1000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted cpu/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module <= cpu_data_master_saved_grant_cpu_jtag_debug_module ? 1 : (cpu_jtag_debug_module_arbitration_holdoff_internal | ~cpu_data_master_requests_cpu_jtag_debug_module) ? 0 : last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module & cpu_data_master_requests_cpu_jtag_debug_module;

  assign cpu_instruction_master_qualified_request_cpu_jtag_debug_module = cpu_instruction_master_requests_cpu_jtag_debug_module & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (|cpu_instruction_master_read_data_valid_sdram_s1_shift_register))) | cpu_data_master_arbiterlock);
  //local readdatavalid cpu_instruction_master_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  assign cpu_instruction_master_read_data_valid_cpu_jtag_debug_module = cpu_instruction_master_granted_cpu_jtag_debug_module & cpu_instruction_master_read & ~cpu_jtag_debug_module_waits_for_read;

  //allow new arb cycle for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock;

  //cpu/instruction_master assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_master_qreq_vector[0] = cpu_instruction_master_qualified_request_cpu_jtag_debug_module;

  //cpu/instruction_master grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_instruction_master_granted_cpu_jtag_debug_module = cpu_jtag_debug_module_grant_vector[0];

  //cpu/instruction_master saved-grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_instruction_master_saved_grant_cpu_jtag_debug_module = cpu_jtag_debug_module_arb_winner[0] && cpu_instruction_master_requests_cpu_jtag_debug_module;

  //cpu/data_master assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_master_qreq_vector[1] = cpu_data_master_qualified_request_cpu_jtag_debug_module;

  //cpu/data_master grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_data_master_granted_cpu_jtag_debug_module = cpu_jtag_debug_module_grant_vector[1];

  //cpu/data_master saved-grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_data_master_saved_grant_cpu_jtag_debug_module = cpu_jtag_debug_module_arb_winner[1] && cpu_data_master_requests_cpu_jtag_debug_module;

  //cpu/jtag_debug_module chosen-master double-vector, which is an e_assign
  assign cpu_jtag_debug_module_chosen_master_double_vector = {cpu_jtag_debug_module_master_qreq_vector, cpu_jtag_debug_module_master_qreq_vector} & ({~cpu_jtag_debug_module_master_qreq_vector, ~cpu_jtag_debug_module_master_qreq_vector} + cpu_jtag_debug_module_arb_addend);

  //stable onehot encoding of arb winner
  assign cpu_jtag_debug_module_arb_winner = (cpu_jtag_debug_module_allow_new_arb_cycle & | cpu_jtag_debug_module_grant_vector) ? cpu_jtag_debug_module_grant_vector : cpu_jtag_debug_module_saved_chosen_master_vector;

  //saved cpu_jtag_debug_module_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_saved_chosen_master_vector <= 0;
      else if (cpu_jtag_debug_module_allow_new_arb_cycle)
          cpu_jtag_debug_module_saved_chosen_master_vector <= |cpu_jtag_debug_module_grant_vector ? cpu_jtag_debug_module_grant_vector : cpu_jtag_debug_module_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign cpu_jtag_debug_module_grant_vector = {(cpu_jtag_debug_module_chosen_master_double_vector[1] | cpu_jtag_debug_module_chosen_master_double_vector[3]),
    (cpu_jtag_debug_module_chosen_master_double_vector[0] | cpu_jtag_debug_module_chosen_master_double_vector[2])};

  //cpu/jtag_debug_module chosen master rotated left, which is an e_assign
  assign cpu_jtag_debug_module_chosen_master_rot_left = (cpu_jtag_debug_module_arb_winner << 1) ? (cpu_jtag_debug_module_arb_winner << 1) : 1;

  //cpu/jtag_debug_module's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_arb_addend <= 1;
      else if (|cpu_jtag_debug_module_grant_vector)
          cpu_jtag_debug_module_arb_addend <= cpu_jtag_debug_module_end_xfer? cpu_jtag_debug_module_chosen_master_rot_left : cpu_jtag_debug_module_grant_vector;
    end


  assign cpu_jtag_debug_module_begintransfer = cpu_jtag_debug_module_begins_xfer;
  //cpu_jtag_debug_module_reset_n assignment, which is an e_assign
  assign cpu_jtag_debug_module_reset_n = reset_n;

  //assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest;

  assign cpu_jtag_debug_module_chipselect = cpu_data_master_granted_cpu_jtag_debug_module | cpu_instruction_master_granted_cpu_jtag_debug_module;
  //cpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_firsttransfer = cpu_jtag_debug_module_begins_xfer ? cpu_jtag_debug_module_unreg_firsttransfer : cpu_jtag_debug_module_reg_firsttransfer;

  //cpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_unreg_firsttransfer = ~(cpu_jtag_debug_module_slavearbiterlockenable & cpu_jtag_debug_module_any_continuerequest);

  //cpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_jtag_debug_module_begins_xfer)
          cpu_jtag_debug_module_reg_firsttransfer <= cpu_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_jtag_debug_module_beginbursttransfer_internal = cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign cpu_jtag_debug_module_arbitration_holdoff_internal = cpu_jtag_debug_module_begins_xfer & cpu_jtag_debug_module_firsttransfer;

  //cpu_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_jtag_debug_module_write = cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_write;

  assign shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master = cpu_data_master_address_to_slave;
  //cpu_jtag_debug_module_address mux, which is an e_mux
  assign cpu_jtag_debug_module_address = (cpu_data_master_granted_cpu_jtag_debug_module)? (shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master >> 2) :
    (shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master >> 2);

  assign shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  //d1_cpu_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_jtag_debug_module_end_xfer <= 1;
      else 
        d1_cpu_jtag_debug_module_end_xfer <= cpu_jtag_debug_module_end_xfer;
    end


  //cpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_read = cpu_jtag_debug_module_in_a_read_cycle & cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_read_cycle = (cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_read) | (cpu_instruction_master_granted_cpu_jtag_debug_module & cpu_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_jtag_debug_module_in_a_read_cycle;

  //cpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_write = cpu_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_write_cycle = cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_jtag_debug_module_counter = 0;
  //cpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_jtag_debug_module_byteenable = (cpu_data_master_granted_cpu_jtag_debug_module)? cpu_data_master_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_jtag_debug_module_debugaccess = (cpu_data_master_granted_cpu_jtag_debug_module)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_cpu_jtag_debug_module + cpu_instruction_master_granted_cpu_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_cpu_jtag_debug_module + cpu_instruction_master_saved_grant_cpu_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_data_master_arbitrator (
                                    // inputs:
                                     PIO_LCD_B_s1_readdata_from_sa,
                                     PIO_LCD_CLK_s1_readdata_from_sa,
                                     PIO_LCD_CTRL_s1_readdata_from_sa,
                                     PIO_LCD_G_s1_readdata_from_sa,
                                     PIO_LCD_PWM_s1_readdata_from_sa,
                                     PIO_LCD_R_s1_readdata_from_sa,
                                     PIO_LED_s1_readdata_from_sa,
                                     RS232_s1_irq_from_sa,
                                     RS232_s1_readdata_from_sa,
                                     clk,
                                     cpu_data_master_address,
                                     cpu_data_master_byteenable_sdram_s1,
                                     cpu_data_master_granted_PIO_LCD_B_s1,
                                     cpu_data_master_granted_PIO_LCD_CLK_s1,
                                     cpu_data_master_granted_PIO_LCD_CTRL_s1,
                                     cpu_data_master_granted_PIO_LCD_G_s1,
                                     cpu_data_master_granted_PIO_LCD_PWM_s1,
                                     cpu_data_master_granted_PIO_LCD_R_s1,
                                     cpu_data_master_granted_PIO_LED_s1,
                                     cpu_data_master_granted_RS232_s1,
                                     cpu_data_master_granted_cpu_jtag_debug_module,
                                     cpu_data_master_granted_epcs_epcs_control_port,
                                     cpu_data_master_granted_jtag_uart_avalon_jtag_slave,
                                     cpu_data_master_granted_sdram_s1,
                                     cpu_data_master_granted_sysid_control_slave,
                                     cpu_data_master_qualified_request_PIO_LCD_B_s1,
                                     cpu_data_master_qualified_request_PIO_LCD_CLK_s1,
                                     cpu_data_master_qualified_request_PIO_LCD_CTRL_s1,
                                     cpu_data_master_qualified_request_PIO_LCD_G_s1,
                                     cpu_data_master_qualified_request_PIO_LCD_PWM_s1,
                                     cpu_data_master_qualified_request_PIO_LCD_R_s1,
                                     cpu_data_master_qualified_request_PIO_LED_s1,
                                     cpu_data_master_qualified_request_RS232_s1,
                                     cpu_data_master_qualified_request_cpu_jtag_debug_module,
                                     cpu_data_master_qualified_request_epcs_epcs_control_port,
                                     cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave,
                                     cpu_data_master_qualified_request_sdram_s1,
                                     cpu_data_master_qualified_request_sysid_control_slave,
                                     cpu_data_master_read,
                                     cpu_data_master_read_data_valid_PIO_LCD_B_s1,
                                     cpu_data_master_read_data_valid_PIO_LCD_CLK_s1,
                                     cpu_data_master_read_data_valid_PIO_LCD_CTRL_s1,
                                     cpu_data_master_read_data_valid_PIO_LCD_G_s1,
                                     cpu_data_master_read_data_valid_PIO_LCD_PWM_s1,
                                     cpu_data_master_read_data_valid_PIO_LCD_R_s1,
                                     cpu_data_master_read_data_valid_PIO_LED_s1,
                                     cpu_data_master_read_data_valid_RS232_s1,
                                     cpu_data_master_read_data_valid_cpu_jtag_debug_module,
                                     cpu_data_master_read_data_valid_epcs_epcs_control_port,
                                     cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave,
                                     cpu_data_master_read_data_valid_sdram_s1,
                                     cpu_data_master_read_data_valid_sdram_s1_shift_register,
                                     cpu_data_master_read_data_valid_sysid_control_slave,
                                     cpu_data_master_requests_PIO_LCD_B_s1,
                                     cpu_data_master_requests_PIO_LCD_CLK_s1,
                                     cpu_data_master_requests_PIO_LCD_CTRL_s1,
                                     cpu_data_master_requests_PIO_LCD_G_s1,
                                     cpu_data_master_requests_PIO_LCD_PWM_s1,
                                     cpu_data_master_requests_PIO_LCD_R_s1,
                                     cpu_data_master_requests_PIO_LED_s1,
                                     cpu_data_master_requests_RS232_s1,
                                     cpu_data_master_requests_cpu_jtag_debug_module,
                                     cpu_data_master_requests_epcs_epcs_control_port,
                                     cpu_data_master_requests_jtag_uart_avalon_jtag_slave,
                                     cpu_data_master_requests_sdram_s1,
                                     cpu_data_master_requests_sysid_control_slave,
                                     cpu_data_master_write,
                                     cpu_data_master_writedata,
                                     cpu_jtag_debug_module_readdata_from_sa,
                                     d1_PIO_LCD_B_s1_end_xfer,
                                     d1_PIO_LCD_CLK_s1_end_xfer,
                                     d1_PIO_LCD_CTRL_s1_end_xfer,
                                     d1_PIO_LCD_G_s1_end_xfer,
                                     d1_PIO_LCD_PWM_s1_end_xfer,
                                     d1_PIO_LCD_R_s1_end_xfer,
                                     d1_PIO_LED_s1_end_xfer,
                                     d1_RS232_s1_end_xfer,
                                     d1_cpu_jtag_debug_module_end_xfer,
                                     d1_epcs_epcs_control_port_end_xfer,
                                     d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                     d1_sdram_s1_end_xfer,
                                     d1_sysid_control_slave_end_xfer,
                                     epcs_epcs_control_port_irq_from_sa,
                                     epcs_epcs_control_port_readdata_from_sa,
                                     jtag_uart_avalon_jtag_slave_irq_from_sa,
                                     jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                     jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                     reset_n,
                                     sdram_s1_readdata_from_sa,
                                     sdram_s1_waitrequest_from_sa,
                                     sysid_control_slave_readdata_from_sa,

                                    // outputs:
                                     cpu_data_master_address_to_slave,
                                     cpu_data_master_dbs_address,
                                     cpu_data_master_dbs_write_16,
                                     cpu_data_master_irq,
                                     cpu_data_master_no_byte_enables_and_last_term,
                                     cpu_data_master_readdata,
                                     cpu_data_master_waitrequest
                                  )
;

  output  [ 26: 0] cpu_data_master_address_to_slave;
  output  [  1: 0] cpu_data_master_dbs_address;
  output  [ 15: 0] cpu_data_master_dbs_write_16;
  output  [ 31: 0] cpu_data_master_irq;
  output           cpu_data_master_no_byte_enables_and_last_term;
  output  [ 31: 0] cpu_data_master_readdata;
  output           cpu_data_master_waitrequest;
  input   [ 31: 0] PIO_LCD_B_s1_readdata_from_sa;
  input   [ 31: 0] PIO_LCD_CLK_s1_readdata_from_sa;
  input   [ 31: 0] PIO_LCD_CTRL_s1_readdata_from_sa;
  input   [ 31: 0] PIO_LCD_G_s1_readdata_from_sa;
  input   [ 31: 0] PIO_LCD_PWM_s1_readdata_from_sa;
  input   [ 31: 0] PIO_LCD_R_s1_readdata_from_sa;
  input   [ 31: 0] PIO_LED_s1_readdata_from_sa;
  input            RS232_s1_irq_from_sa;
  input   [ 15: 0] RS232_s1_readdata_from_sa;
  input            clk;
  input   [ 26: 0] cpu_data_master_address;
  input   [  1: 0] cpu_data_master_byteenable_sdram_s1;
  input            cpu_data_master_granted_PIO_LCD_B_s1;
  input            cpu_data_master_granted_PIO_LCD_CLK_s1;
  input            cpu_data_master_granted_PIO_LCD_CTRL_s1;
  input            cpu_data_master_granted_PIO_LCD_G_s1;
  input            cpu_data_master_granted_PIO_LCD_PWM_s1;
  input            cpu_data_master_granted_PIO_LCD_R_s1;
  input            cpu_data_master_granted_PIO_LED_s1;
  input            cpu_data_master_granted_RS232_s1;
  input            cpu_data_master_granted_cpu_jtag_debug_module;
  input            cpu_data_master_granted_epcs_epcs_control_port;
  input            cpu_data_master_granted_jtag_uart_avalon_jtag_slave;
  input            cpu_data_master_granted_sdram_s1;
  input            cpu_data_master_granted_sysid_control_slave;
  input            cpu_data_master_qualified_request_PIO_LCD_B_s1;
  input            cpu_data_master_qualified_request_PIO_LCD_CLK_s1;
  input            cpu_data_master_qualified_request_PIO_LCD_CTRL_s1;
  input            cpu_data_master_qualified_request_PIO_LCD_G_s1;
  input            cpu_data_master_qualified_request_PIO_LCD_PWM_s1;
  input            cpu_data_master_qualified_request_PIO_LCD_R_s1;
  input            cpu_data_master_qualified_request_PIO_LED_s1;
  input            cpu_data_master_qualified_request_RS232_s1;
  input            cpu_data_master_qualified_request_cpu_jtag_debug_module;
  input            cpu_data_master_qualified_request_epcs_epcs_control_port;
  input            cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave;
  input            cpu_data_master_qualified_request_sdram_s1;
  input            cpu_data_master_qualified_request_sysid_control_slave;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_PIO_LCD_B_s1;
  input            cpu_data_master_read_data_valid_PIO_LCD_CLK_s1;
  input            cpu_data_master_read_data_valid_PIO_LCD_CTRL_s1;
  input            cpu_data_master_read_data_valid_PIO_LCD_G_s1;
  input            cpu_data_master_read_data_valid_PIO_LCD_PWM_s1;
  input            cpu_data_master_read_data_valid_PIO_LCD_R_s1;
  input            cpu_data_master_read_data_valid_PIO_LED_s1;
  input            cpu_data_master_read_data_valid_RS232_s1;
  input            cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  input            cpu_data_master_read_data_valid_epcs_epcs_control_port;
  input            cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave;
  input            cpu_data_master_read_data_valid_sdram_s1;
  input            cpu_data_master_read_data_valid_sdram_s1_shift_register;
  input            cpu_data_master_read_data_valid_sysid_control_slave;
  input            cpu_data_master_requests_PIO_LCD_B_s1;
  input            cpu_data_master_requests_PIO_LCD_CLK_s1;
  input            cpu_data_master_requests_PIO_LCD_CTRL_s1;
  input            cpu_data_master_requests_PIO_LCD_G_s1;
  input            cpu_data_master_requests_PIO_LCD_PWM_s1;
  input            cpu_data_master_requests_PIO_LCD_R_s1;
  input            cpu_data_master_requests_PIO_LED_s1;
  input            cpu_data_master_requests_RS232_s1;
  input            cpu_data_master_requests_cpu_jtag_debug_module;
  input            cpu_data_master_requests_epcs_epcs_control_port;
  input            cpu_data_master_requests_jtag_uart_avalon_jtag_slave;
  input            cpu_data_master_requests_sdram_s1;
  input            cpu_data_master_requests_sysid_control_slave;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  input            d1_PIO_LCD_B_s1_end_xfer;
  input            d1_PIO_LCD_CLK_s1_end_xfer;
  input            d1_PIO_LCD_CTRL_s1_end_xfer;
  input            d1_PIO_LCD_G_s1_end_xfer;
  input            d1_PIO_LCD_PWM_s1_end_xfer;
  input            d1_PIO_LCD_R_s1_end_xfer;
  input            d1_PIO_LED_s1_end_xfer;
  input            d1_RS232_s1_end_xfer;
  input            d1_cpu_jtag_debug_module_end_xfer;
  input            d1_epcs_epcs_control_port_end_xfer;
  input            d1_jtag_uart_avalon_jtag_slave_end_xfer;
  input            d1_sdram_s1_end_xfer;
  input            d1_sysid_control_slave_end_xfer;
  input            epcs_epcs_control_port_irq_from_sa;
  input   [ 31: 0] epcs_epcs_control_port_readdata_from_sa;
  input            jtag_uart_avalon_jtag_slave_irq_from_sa;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  input            reset_n;
  input   [ 15: 0] sdram_s1_readdata_from_sa;
  input            sdram_s1_waitrequest_from_sa;
  input   [ 31: 0] sysid_control_slave_readdata_from_sa;

  wire    [ 26: 0] cpu_data_master_address_to_slave;
  reg     [  1: 0] cpu_data_master_dbs_address;
  wire    [  1: 0] cpu_data_master_dbs_increment;
  wire    [ 15: 0] cpu_data_master_dbs_write_16;
  wire    [ 31: 0] cpu_data_master_irq;
  reg              cpu_data_master_no_byte_enables_and_last_term;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_run;
  reg              cpu_data_master_waitrequest;
  reg     [ 15: 0] dbs_16_reg_segment_0;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  wire             last_dbs_term_and_run;
  wire    [  1: 0] next_dbs_address;
  wire    [ 15: 0] p1_dbs_16_reg_segment_0;
  wire    [ 31: 0] p1_registered_cpu_data_master_readdata;
  wire             pre_dbs_count_enable;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  reg     [ 31: 0] registered_cpu_data_master_readdata;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_data_master_qualified_request_PIO_LCD_B_s1 | ~cpu_data_master_requests_PIO_LCD_B_s1) & ((~cpu_data_master_qualified_request_PIO_LCD_B_s1 | ~cpu_data_master_read | (1 & 1 & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_PIO_LCD_B_s1 | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_PIO_LCD_CLK_s1 | ~cpu_data_master_requests_PIO_LCD_CLK_s1) & ((~cpu_data_master_qualified_request_PIO_LCD_CLK_s1 | ~cpu_data_master_read | (1 & 1 & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_PIO_LCD_CLK_s1 | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_PIO_LCD_CTRL_s1 | ~cpu_data_master_requests_PIO_LCD_CTRL_s1) & ((~cpu_data_master_qualified_request_PIO_LCD_CTRL_s1 | ~cpu_data_master_read | (1 & 1 & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_PIO_LCD_CTRL_s1 | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_PIO_LCD_G_s1 | ~cpu_data_master_requests_PIO_LCD_G_s1) & ((~cpu_data_master_qualified_request_PIO_LCD_G_s1 | ~cpu_data_master_read | (1 & 1 & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_PIO_LCD_G_s1 | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_PIO_LCD_PWM_s1 | ~cpu_data_master_requests_PIO_LCD_PWM_s1) & ((~cpu_data_master_qualified_request_PIO_LCD_PWM_s1 | ~cpu_data_master_read | (1 & 1 & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_PIO_LCD_PWM_s1 | ~cpu_data_master_write | (1 & cpu_data_master_write)));

  //cascaded wait assignment, which is an e_assign
  assign cpu_data_master_run = r_0 & r_1 & r_2;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_data_master_qualified_request_PIO_LCD_R_s1 | ~cpu_data_master_requests_PIO_LCD_R_s1) & ((~cpu_data_master_qualified_request_PIO_LCD_R_s1 | ~cpu_data_master_read | (1 & 1 & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_PIO_LCD_R_s1 | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_PIO_LED_s1 | ~cpu_data_master_requests_PIO_LED_s1) & ((~cpu_data_master_qualified_request_PIO_LED_s1 | ~cpu_data_master_read | (1 & 1 & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_PIO_LED_s1 | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & ((~cpu_data_master_qualified_request_RS232_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & 1 & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_RS232_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & 1 & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_cpu_jtag_debug_module | ~cpu_data_master_requests_cpu_jtag_debug_module) & (cpu_data_master_granted_cpu_jtag_debug_module | ~cpu_data_master_qualified_request_cpu_jtag_debug_module) & ((~cpu_data_master_qualified_request_cpu_jtag_debug_module | ~cpu_data_master_read | (1 & 1 & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_cpu_jtag_debug_module | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_epcs_epcs_control_port | ~cpu_data_master_requests_epcs_epcs_control_port) & (cpu_data_master_granted_epcs_epcs_control_port | ~cpu_data_master_qualified_request_epcs_epcs_control_port) & ((~cpu_data_master_qualified_request_epcs_epcs_control_port | ~(cpu_data_master_read | cpu_data_master_write) | (1 & 1 & (cpu_data_master_read | cpu_data_master_write))));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = ((~cpu_data_master_qualified_request_epcs_epcs_control_port | ~(cpu_data_master_read | cpu_data_master_write) | (1 & 1 & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave | ~cpu_data_master_requests_jtag_uart_avalon_jtag_slave) & ((~cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_sdram_s1 | (cpu_data_master_read_data_valid_sdram_s1 & cpu_data_master_dbs_address[1]) | (cpu_data_master_write & !cpu_data_master_byteenable_sdram_s1 & cpu_data_master_dbs_address[1]) | ~cpu_data_master_requests_sdram_s1) & (cpu_data_master_granted_sdram_s1 | ~cpu_data_master_qualified_request_sdram_s1) & ((~cpu_data_master_qualified_request_sdram_s1 | ~cpu_data_master_read | (cpu_data_master_read_data_valid_sdram_s1 & (cpu_data_master_dbs_address[1]) & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_sdram_s1 | ~cpu_data_master_write | (1 & ~sdram_s1_waitrequest_from_sa & (cpu_data_master_dbs_address[1]) & cpu_data_master_write))) & 1 & ((~cpu_data_master_qualified_request_sysid_control_slave | ~cpu_data_master_read | (1 & 1 & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_sysid_control_slave | ~cpu_data_master_write | (1 & cpu_data_master_write)));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_data_master_address_to_slave = {cpu_data_master_address[26],
    1'b0,
    cpu_data_master_address[24 : 0]};

  //cpu/data_master readdata mux, which is an e_mux
  assign cpu_data_master_readdata = ({32 {~cpu_data_master_requests_PIO_LCD_B_s1}} | PIO_LCD_B_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_requests_PIO_LCD_CLK_s1}} | PIO_LCD_CLK_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_requests_PIO_LCD_CTRL_s1}} | PIO_LCD_CTRL_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_requests_PIO_LCD_G_s1}} | PIO_LCD_G_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_requests_PIO_LCD_PWM_s1}} | PIO_LCD_PWM_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_requests_PIO_LCD_R_s1}} | PIO_LCD_R_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_requests_PIO_LED_s1}} | PIO_LED_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_requests_RS232_s1}} | RS232_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_requests_cpu_jtag_debug_module}} | cpu_jtag_debug_module_readdata_from_sa) &
    ({32 {~cpu_data_master_requests_epcs_epcs_control_port}} | epcs_epcs_control_port_readdata_from_sa) &
    ({32 {~cpu_data_master_requests_jtag_uart_avalon_jtag_slave}} | registered_cpu_data_master_readdata) &
    ({32 {~cpu_data_master_requests_sdram_s1}} | registered_cpu_data_master_readdata) &
    ({32 {~cpu_data_master_requests_sysid_control_slave}} | sysid_control_slave_readdata_from_sa);

  //actual waitrequest port, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_waitrequest <= ~0;
      else 
        cpu_data_master_waitrequest <= ~((~(cpu_data_master_read | cpu_data_master_write))? 0: (cpu_data_master_run & cpu_data_master_waitrequest));
    end


  //irq assign, which is an e_assign
  assign cpu_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    RS232_s1_irq_from_sa,
    jtag_uart_avalon_jtag_slave_irq_from_sa,
    epcs_epcs_control_port_irq_from_sa};

  //unpredictable registered wait state incoming data, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_cpu_data_master_readdata <= 0;
      else 
        registered_cpu_data_master_readdata <= p1_registered_cpu_data_master_readdata;
    end


  //registered readdata mux, which is an e_mux
  assign p1_registered_cpu_data_master_readdata = ({32 {~cpu_data_master_requests_jtag_uart_avalon_jtag_slave}} | jtag_uart_avalon_jtag_slave_readdata_from_sa) &
    ({32 {~cpu_data_master_requests_sdram_s1}} | {sdram_s1_readdata_from_sa[15 : 0],
    dbs_16_reg_segment_0});

  //no_byte_enables_and_last_term, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_no_byte_enables_and_last_term <= 0;
      else 
        cpu_data_master_no_byte_enables_and_last_term <= last_dbs_term_and_run;
    end


  //compute the last dbs term, which is an e_mux
  assign last_dbs_term_and_run = (cpu_data_master_dbs_address == 2'b10) & cpu_data_master_write & !cpu_data_master_byteenable_sdram_s1;

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (((~cpu_data_master_no_byte_enables_and_last_term) & cpu_data_master_requests_sdram_s1 & cpu_data_master_write & !cpu_data_master_byteenable_sdram_s1)) |
    cpu_data_master_read_data_valid_sdram_s1 |
    (cpu_data_master_granted_sdram_s1 & cpu_data_master_write & 1 & 1 & ~sdram_s1_waitrequest_from_sa);

  //input to dbs-16 stored 0, which is an e_mux
  assign p1_dbs_16_reg_segment_0 = sdram_s1_readdata_from_sa;

  //dbs register for dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_16_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_data_master_dbs_address[1]) == 0))
          dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
    end


  //mux write dbs 1, which is an e_mux
  assign cpu_data_master_dbs_write_16 = (cpu_data_master_dbs_address[1])? cpu_data_master_writedata[31 : 16] :
    cpu_data_master_writedata[15 : 0];

  //dbs count increment, which is an e_mux
  assign cpu_data_master_dbs_increment = (cpu_data_master_requests_sdram_s1)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_data_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_data_master_dbs_address + cpu_data_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable &
    (~(cpu_data_master_requests_sdram_s1 & ~cpu_data_master_waitrequest));

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_data_master_dbs_address <= next_dbs_address;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_instruction_master_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_instruction_master_address,
                                            cpu_instruction_master_granted_cpu_jtag_debug_module,
                                            cpu_instruction_master_granted_epcs_epcs_control_port,
                                            cpu_instruction_master_granted_sdram_s1,
                                            cpu_instruction_master_qualified_request_cpu_jtag_debug_module,
                                            cpu_instruction_master_qualified_request_epcs_epcs_control_port,
                                            cpu_instruction_master_qualified_request_sdram_s1,
                                            cpu_instruction_master_read,
                                            cpu_instruction_master_read_data_valid_cpu_jtag_debug_module,
                                            cpu_instruction_master_read_data_valid_epcs_epcs_control_port,
                                            cpu_instruction_master_read_data_valid_sdram_s1,
                                            cpu_instruction_master_read_data_valid_sdram_s1_shift_register,
                                            cpu_instruction_master_requests_cpu_jtag_debug_module,
                                            cpu_instruction_master_requests_epcs_epcs_control_port,
                                            cpu_instruction_master_requests_sdram_s1,
                                            cpu_jtag_debug_module_readdata_from_sa,
                                            d1_cpu_jtag_debug_module_end_xfer,
                                            d1_epcs_epcs_control_port_end_xfer,
                                            d1_sdram_s1_end_xfer,
                                            epcs_epcs_control_port_readdata_from_sa,
                                            reset_n,
                                            sdram_s1_readdata_from_sa,
                                            sdram_s1_waitrequest_from_sa,

                                           // outputs:
                                            cpu_instruction_master_address_to_slave,
                                            cpu_instruction_master_dbs_address,
                                            cpu_instruction_master_latency_counter,
                                            cpu_instruction_master_readdata,
                                            cpu_instruction_master_readdatavalid,
                                            cpu_instruction_master_waitrequest
                                         )
;

  output  [ 26: 0] cpu_instruction_master_address_to_slave;
  output  [  1: 0] cpu_instruction_master_dbs_address;
  output           cpu_instruction_master_latency_counter;
  output  [ 31: 0] cpu_instruction_master_readdata;
  output           cpu_instruction_master_readdatavalid;
  output           cpu_instruction_master_waitrequest;
  input            clk;
  input   [ 26: 0] cpu_instruction_master_address;
  input            cpu_instruction_master_granted_cpu_jtag_debug_module;
  input            cpu_instruction_master_granted_epcs_epcs_control_port;
  input            cpu_instruction_master_granted_sdram_s1;
  input            cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  input            cpu_instruction_master_qualified_request_epcs_epcs_control_port;
  input            cpu_instruction_master_qualified_request_sdram_s1;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  input            cpu_instruction_master_read_data_valid_epcs_epcs_control_port;
  input            cpu_instruction_master_read_data_valid_sdram_s1;
  input            cpu_instruction_master_read_data_valid_sdram_s1_shift_register;
  input            cpu_instruction_master_requests_cpu_jtag_debug_module;
  input            cpu_instruction_master_requests_epcs_epcs_control_port;
  input            cpu_instruction_master_requests_sdram_s1;
  input   [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_jtag_debug_module_end_xfer;
  input            d1_epcs_epcs_control_port_end_xfer;
  input            d1_sdram_s1_end_xfer;
  input   [ 31: 0] epcs_epcs_control_port_readdata_from_sa;
  input            reset_n;
  input   [ 15: 0] sdram_s1_readdata_from_sa;
  input            sdram_s1_waitrequest_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 26: 0] cpu_instruction_master_address_last_time;
  wire    [ 26: 0] cpu_instruction_master_address_to_slave;
  reg     [  1: 0] cpu_instruction_master_dbs_address;
  wire    [  1: 0] cpu_instruction_master_dbs_increment;
  reg     [  1: 0] cpu_instruction_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_instruction_master_dbs_rdv_counter_inc;
  wire             cpu_instruction_master_is_granted_some_slave;
  reg              cpu_instruction_master_latency_counter;
  wire    [  1: 0] cpu_instruction_master_next_dbs_rdv_counter;
  reg              cpu_instruction_master_read_but_no_slave_selected;
  reg              cpu_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_run;
  wire             cpu_instruction_master_waitrequest;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire             latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire             p1_cpu_instruction_master_latency_counter;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_instruction_master_readdatavalid;
  wire             r_1;
  wire             r_2;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_instruction_master_qualified_request_cpu_jtag_debug_module | ~cpu_instruction_master_requests_cpu_jtag_debug_module) & (cpu_instruction_master_granted_cpu_jtag_debug_module | ~cpu_instruction_master_qualified_request_cpu_jtag_debug_module) & ((~cpu_instruction_master_qualified_request_cpu_jtag_debug_module | ~cpu_instruction_master_read | (1 & ~d1_cpu_jtag_debug_module_end_xfer & cpu_instruction_master_read))) & 1 & (cpu_instruction_master_qualified_request_epcs_epcs_control_port | ~cpu_instruction_master_requests_epcs_epcs_control_port) & (cpu_instruction_master_granted_epcs_epcs_control_port | ~cpu_instruction_master_qualified_request_epcs_epcs_control_port);

  //cascaded wait assignment, which is an e_assign
  assign cpu_instruction_master_run = r_1 & r_2;

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = ((~cpu_instruction_master_qualified_request_epcs_epcs_control_port | ~(cpu_instruction_master_read) | (1 & ~d1_epcs_epcs_control_port_end_xfer & (cpu_instruction_master_read)))) & 1 & (cpu_instruction_master_qualified_request_sdram_s1 | ~cpu_instruction_master_requests_sdram_s1) & (cpu_instruction_master_granted_sdram_s1 | ~cpu_instruction_master_qualified_request_sdram_s1) & ((~cpu_instruction_master_qualified_request_sdram_s1 | ~cpu_instruction_master_read | (1 & ~sdram_s1_waitrequest_from_sa & (cpu_instruction_master_dbs_address[1]) & cpu_instruction_master_read)));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_instruction_master_address_to_slave = {cpu_instruction_master_address[26],
    1'b0,
    cpu_instruction_master_address[24 : 0]};

  //cpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_but_no_slave_selected <= 0;
      else 
        cpu_instruction_master_read_but_no_slave_selected <= cpu_instruction_master_read & cpu_instruction_master_run & ~cpu_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_instruction_master_is_granted_some_slave = cpu_instruction_master_granted_cpu_jtag_debug_module |
    cpu_instruction_master_granted_epcs_epcs_control_port |
    cpu_instruction_master_granted_sdram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_instruction_master_readdatavalid = cpu_instruction_master_read_data_valid_sdram_s1 & dbs_rdv_counter_overflow;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_instruction_master_readdatavalid = cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_data_valid_cpu_jtag_debug_module |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_data_valid_epcs_epcs_control_port |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid;

  //cpu/instruction_master readdata mux, which is an e_mux
  assign cpu_instruction_master_readdata = ({32 {~(cpu_instruction_master_qualified_request_cpu_jtag_debug_module & cpu_instruction_master_read)}} | cpu_jtag_debug_module_readdata_from_sa) &
    ({32 {~(cpu_instruction_master_qualified_request_epcs_epcs_control_port & cpu_instruction_master_read)}} | epcs_epcs_control_port_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_sdram_s1}} | {sdram_s1_readdata_from_sa[15 : 0],
    dbs_latent_16_reg_segment_0});

  //actual waitrequest port, which is an e_assign
  assign cpu_instruction_master_waitrequest = ~cpu_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_latency_counter <= 0;
      else 
        cpu_instruction_master_latency_counter <= p1_cpu_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_instruction_master_latency_counter = ((cpu_instruction_master_run & cpu_instruction_master_read))? latency_load_value :
    (cpu_instruction_master_latency_counter)? cpu_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = sdram_s1_readdata_from_sa;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_instruction_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //dbs count increment, which is an e_mux
  assign cpu_instruction_master_dbs_increment = (cpu_instruction_master_requests_sdram_s1)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_instruction_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_instruction_master_dbs_address + cpu_instruction_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_instruction_master_dbs_address <= next_dbs_address;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_instruction_master_next_dbs_rdv_counter = cpu_instruction_master_dbs_rdv_counter + cpu_instruction_master_dbs_rdv_counter_inc;

  //cpu_instruction_master_rdv_inc_mux, which is an e_mux
  assign cpu_instruction_master_dbs_rdv_counter_inc = 2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_instruction_master_read_data_valid_sdram_s1;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_instruction_master_dbs_rdv_counter <= cpu_instruction_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_instruction_master_dbs_rdv_counter[1] & ~cpu_instruction_master_next_dbs_rdv_counter[1];

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = cpu_instruction_master_granted_sdram_s1 & cpu_instruction_master_read & 1 & 1 & ~sdram_s1_waitrequest_from_sa;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_address_last_time <= 0;
      else 
        cpu_instruction_master_address_last_time <= cpu_instruction_master_address;
    end


  //cpu/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_instruction_master_waitrequest & (cpu_instruction_master_read);
    end


  //cpu_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_address != cpu_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_last_time <= 0;
      else 
        cpu_instruction_master_read_last_time <= cpu_instruction_master_read;
    end


  //cpu_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_read != cpu_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module epcs_epcs_control_port_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_data_master_address_to_slave,
                                            cpu_data_master_read,
                                            cpu_data_master_write,
                                            cpu_data_master_writedata,
                                            cpu_instruction_master_address_to_slave,
                                            cpu_instruction_master_latency_counter,
                                            cpu_instruction_master_read,
                                            cpu_instruction_master_read_data_valid_sdram_s1_shift_register,
                                            epcs_epcs_control_port_dataavailable,
                                            epcs_epcs_control_port_endofpacket,
                                            epcs_epcs_control_port_irq,
                                            epcs_epcs_control_port_readdata,
                                            epcs_epcs_control_port_readyfordata,
                                            reset_n,

                                           // outputs:
                                            cpu_data_master_granted_epcs_epcs_control_port,
                                            cpu_data_master_qualified_request_epcs_epcs_control_port,
                                            cpu_data_master_read_data_valid_epcs_epcs_control_port,
                                            cpu_data_master_requests_epcs_epcs_control_port,
                                            cpu_instruction_master_granted_epcs_epcs_control_port,
                                            cpu_instruction_master_qualified_request_epcs_epcs_control_port,
                                            cpu_instruction_master_read_data_valid_epcs_epcs_control_port,
                                            cpu_instruction_master_requests_epcs_epcs_control_port,
                                            d1_epcs_epcs_control_port_end_xfer,
                                            epcs_epcs_control_port_address,
                                            epcs_epcs_control_port_chipselect,
                                            epcs_epcs_control_port_dataavailable_from_sa,
                                            epcs_epcs_control_port_endofpacket_from_sa,
                                            epcs_epcs_control_port_irq_from_sa,
                                            epcs_epcs_control_port_read_n,
                                            epcs_epcs_control_port_readdata_from_sa,
                                            epcs_epcs_control_port_readyfordata_from_sa,
                                            epcs_epcs_control_port_reset_n,
                                            epcs_epcs_control_port_write_n,
                                            epcs_epcs_control_port_writedata
                                         )
;

  output           cpu_data_master_granted_epcs_epcs_control_port;
  output           cpu_data_master_qualified_request_epcs_epcs_control_port;
  output           cpu_data_master_read_data_valid_epcs_epcs_control_port;
  output           cpu_data_master_requests_epcs_epcs_control_port;
  output           cpu_instruction_master_granted_epcs_epcs_control_port;
  output           cpu_instruction_master_qualified_request_epcs_epcs_control_port;
  output           cpu_instruction_master_read_data_valid_epcs_epcs_control_port;
  output           cpu_instruction_master_requests_epcs_epcs_control_port;
  output           d1_epcs_epcs_control_port_end_xfer;
  output  [  8: 0] epcs_epcs_control_port_address;
  output           epcs_epcs_control_port_chipselect;
  output           epcs_epcs_control_port_dataavailable_from_sa;
  output           epcs_epcs_control_port_endofpacket_from_sa;
  output           epcs_epcs_control_port_irq_from_sa;
  output           epcs_epcs_control_port_read_n;
  output  [ 31: 0] epcs_epcs_control_port_readdata_from_sa;
  output           epcs_epcs_control_port_readyfordata_from_sa;
  output           epcs_epcs_control_port_reset_n;
  output           epcs_epcs_control_port_write_n;
  output  [ 31: 0] epcs_epcs_control_port_writedata;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_read;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 26: 0] cpu_instruction_master_address_to_slave;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_sdram_s1_shift_register;
  input            epcs_epcs_control_port_dataavailable;
  input            epcs_epcs_control_port_endofpacket;
  input            epcs_epcs_control_port_irq;
  input   [ 31: 0] epcs_epcs_control_port_readdata;
  input            epcs_epcs_control_port_readyfordata;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_epcs_epcs_control_port;
  wire             cpu_data_master_qualified_request_epcs_epcs_control_port;
  wire             cpu_data_master_read_data_valid_epcs_epcs_control_port;
  wire             cpu_data_master_requests_epcs_epcs_control_port;
  wire             cpu_data_master_saved_grant_epcs_epcs_control_port;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_epcs_epcs_control_port;
  wire             cpu_instruction_master_qualified_request_epcs_epcs_control_port;
  wire             cpu_instruction_master_read_data_valid_epcs_epcs_control_port;
  wire             cpu_instruction_master_requests_epcs_epcs_control_port;
  wire             cpu_instruction_master_saved_grant_epcs_epcs_control_port;
  reg              d1_epcs_epcs_control_port_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_epcs_epcs_control_port;
  wire    [  8: 0] epcs_epcs_control_port_address;
  wire             epcs_epcs_control_port_allgrants;
  wire             epcs_epcs_control_port_allow_new_arb_cycle;
  wire             epcs_epcs_control_port_any_bursting_master_saved_grant;
  wire             epcs_epcs_control_port_any_continuerequest;
  reg     [  1: 0] epcs_epcs_control_port_arb_addend;
  wire             epcs_epcs_control_port_arb_counter_enable;
  reg     [  1: 0] epcs_epcs_control_port_arb_share_counter;
  wire    [  1: 0] epcs_epcs_control_port_arb_share_counter_next_value;
  wire    [  1: 0] epcs_epcs_control_port_arb_share_set_values;
  wire    [  1: 0] epcs_epcs_control_port_arb_winner;
  wire             epcs_epcs_control_port_arbitration_holdoff_internal;
  wire             epcs_epcs_control_port_beginbursttransfer_internal;
  wire             epcs_epcs_control_port_begins_xfer;
  wire             epcs_epcs_control_port_chipselect;
  wire    [  3: 0] epcs_epcs_control_port_chosen_master_double_vector;
  wire    [  1: 0] epcs_epcs_control_port_chosen_master_rot_left;
  wire             epcs_epcs_control_port_dataavailable_from_sa;
  wire             epcs_epcs_control_port_end_xfer;
  wire             epcs_epcs_control_port_endofpacket_from_sa;
  wire             epcs_epcs_control_port_firsttransfer;
  wire    [  1: 0] epcs_epcs_control_port_grant_vector;
  wire             epcs_epcs_control_port_in_a_read_cycle;
  wire             epcs_epcs_control_port_in_a_write_cycle;
  wire             epcs_epcs_control_port_irq_from_sa;
  wire    [  1: 0] epcs_epcs_control_port_master_qreq_vector;
  wire             epcs_epcs_control_port_non_bursting_master_requests;
  wire             epcs_epcs_control_port_read_n;
  wire    [ 31: 0] epcs_epcs_control_port_readdata_from_sa;
  wire             epcs_epcs_control_port_readyfordata_from_sa;
  reg              epcs_epcs_control_port_reg_firsttransfer;
  wire             epcs_epcs_control_port_reset_n;
  reg     [  1: 0] epcs_epcs_control_port_saved_chosen_master_vector;
  reg              epcs_epcs_control_port_slavearbiterlockenable;
  wire             epcs_epcs_control_port_slavearbiterlockenable2;
  wire             epcs_epcs_control_port_unreg_firsttransfer;
  wire             epcs_epcs_control_port_waits_for_read;
  wire             epcs_epcs_control_port_waits_for_write;
  wire             epcs_epcs_control_port_write_n;
  wire    [ 31: 0] epcs_epcs_control_port_writedata;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_epcs_epcs_control_port;
  reg              last_cycle_cpu_instruction_master_granted_slave_epcs_epcs_control_port;
  wire    [ 26: 0] shifted_address_to_epcs_epcs_control_port_from_cpu_data_master;
  wire    [ 26: 0] shifted_address_to_epcs_epcs_control_port_from_cpu_instruction_master;
  wire             wait_for_epcs_epcs_control_port_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~epcs_epcs_control_port_end_xfer;
    end


  assign epcs_epcs_control_port_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_epcs_epcs_control_port | cpu_instruction_master_qualified_request_epcs_epcs_control_port));
  //assign epcs_epcs_control_port_readdata_from_sa = epcs_epcs_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign epcs_epcs_control_port_readdata_from_sa = epcs_epcs_control_port_readdata;

  assign cpu_data_master_requests_epcs_epcs_control_port = ({cpu_data_master_address_to_slave[26 : 11] , 11'b0} == 27'h0) & (cpu_data_master_read | cpu_data_master_write);
  //assign epcs_epcs_control_port_dataavailable_from_sa = epcs_epcs_control_port_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign epcs_epcs_control_port_dataavailable_from_sa = epcs_epcs_control_port_dataavailable;

  //assign epcs_epcs_control_port_readyfordata_from_sa = epcs_epcs_control_port_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign epcs_epcs_control_port_readyfordata_from_sa = epcs_epcs_control_port_readyfordata;

  //epcs_epcs_control_port_arb_share_counter set values, which is an e_mux
  assign epcs_epcs_control_port_arb_share_set_values = 1;

  //epcs_epcs_control_port_non_bursting_master_requests mux, which is an e_mux
  assign epcs_epcs_control_port_non_bursting_master_requests = cpu_data_master_requests_epcs_epcs_control_port |
    cpu_instruction_master_requests_epcs_epcs_control_port |
    cpu_data_master_requests_epcs_epcs_control_port |
    cpu_instruction_master_requests_epcs_epcs_control_port;

  //epcs_epcs_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  assign epcs_epcs_control_port_any_bursting_master_saved_grant = 0;

  //epcs_epcs_control_port_arb_share_counter_next_value assignment, which is an e_assign
  assign epcs_epcs_control_port_arb_share_counter_next_value = epcs_epcs_control_port_firsttransfer ? (epcs_epcs_control_port_arb_share_set_values - 1) : |epcs_epcs_control_port_arb_share_counter ? (epcs_epcs_control_port_arb_share_counter - 1) : 0;

  //epcs_epcs_control_port_allgrants all slave grants, which is an e_mux
  assign epcs_epcs_control_port_allgrants = (|epcs_epcs_control_port_grant_vector) |
    (|epcs_epcs_control_port_grant_vector) |
    (|epcs_epcs_control_port_grant_vector) |
    (|epcs_epcs_control_port_grant_vector);

  //epcs_epcs_control_port_end_xfer assignment, which is an e_assign
  assign epcs_epcs_control_port_end_xfer = ~(epcs_epcs_control_port_waits_for_read | epcs_epcs_control_port_waits_for_write);

  //end_xfer_arb_share_counter_term_epcs_epcs_control_port arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_epcs_epcs_control_port = epcs_epcs_control_port_end_xfer & (~epcs_epcs_control_port_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //epcs_epcs_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  assign epcs_epcs_control_port_arb_counter_enable = (end_xfer_arb_share_counter_term_epcs_epcs_control_port & epcs_epcs_control_port_allgrants) | (end_xfer_arb_share_counter_term_epcs_epcs_control_port & ~epcs_epcs_control_port_non_bursting_master_requests);

  //epcs_epcs_control_port_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          epcs_epcs_control_port_arb_share_counter <= 0;
      else if (epcs_epcs_control_port_arb_counter_enable)
          epcs_epcs_control_port_arb_share_counter <= epcs_epcs_control_port_arb_share_counter_next_value;
    end


  //epcs_epcs_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          epcs_epcs_control_port_slavearbiterlockenable <= 0;
      else if ((|epcs_epcs_control_port_master_qreq_vector & end_xfer_arb_share_counter_term_epcs_epcs_control_port) | (end_xfer_arb_share_counter_term_epcs_epcs_control_port & ~epcs_epcs_control_port_non_bursting_master_requests))
          epcs_epcs_control_port_slavearbiterlockenable <= |epcs_epcs_control_port_arb_share_counter_next_value;
    end


  //cpu/data_master epcs/epcs_control_port arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = epcs_epcs_control_port_slavearbiterlockenable & cpu_data_master_continuerequest;

  //epcs_epcs_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign epcs_epcs_control_port_slavearbiterlockenable2 = |epcs_epcs_control_port_arb_share_counter_next_value;

  //cpu/data_master epcs/epcs_control_port arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = epcs_epcs_control_port_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master epcs/epcs_control_port arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = epcs_epcs_control_port_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master epcs/epcs_control_port arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = epcs_epcs_control_port_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted epcs/epcs_control_port last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_epcs_epcs_control_port <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_epcs_epcs_control_port <= cpu_instruction_master_saved_grant_epcs_epcs_control_port ? 1 : (epcs_epcs_control_port_arbitration_holdoff_internal | ~cpu_instruction_master_requests_epcs_epcs_control_port) ? 0 : last_cycle_cpu_instruction_master_granted_slave_epcs_epcs_control_port;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = last_cycle_cpu_instruction_master_granted_slave_epcs_epcs_control_port & cpu_instruction_master_requests_epcs_epcs_control_port;

  //epcs_epcs_control_port_any_continuerequest at least one master continues requesting, which is an e_mux
  assign epcs_epcs_control_port_any_continuerequest = cpu_instruction_master_continuerequest |
    cpu_data_master_continuerequest;

  assign cpu_data_master_qualified_request_epcs_epcs_control_port = cpu_data_master_requests_epcs_epcs_control_port & ~(cpu_instruction_master_arbiterlock);
  //epcs_epcs_control_port_writedata mux, which is an e_mux
  assign epcs_epcs_control_port_writedata = cpu_data_master_writedata;

  //assign epcs_epcs_control_port_endofpacket_from_sa = epcs_epcs_control_port_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign epcs_epcs_control_port_endofpacket_from_sa = epcs_epcs_control_port_endofpacket;

  assign cpu_instruction_master_requests_epcs_epcs_control_port = (({cpu_instruction_master_address_to_slave[26 : 11] , 11'b0} == 27'h0) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted epcs/epcs_control_port last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_epcs_epcs_control_port <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_epcs_epcs_control_port <= cpu_data_master_saved_grant_epcs_epcs_control_port ? 1 : (epcs_epcs_control_port_arbitration_holdoff_internal | ~cpu_data_master_requests_epcs_epcs_control_port) ? 0 : last_cycle_cpu_data_master_granted_slave_epcs_epcs_control_port;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = last_cycle_cpu_data_master_granted_slave_epcs_epcs_control_port & cpu_data_master_requests_epcs_epcs_control_port;

  assign cpu_instruction_master_qualified_request_epcs_epcs_control_port = cpu_instruction_master_requests_epcs_epcs_control_port & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (|cpu_instruction_master_read_data_valid_sdram_s1_shift_register))) | cpu_data_master_arbiterlock);
  //local readdatavalid cpu_instruction_master_read_data_valid_epcs_epcs_control_port, which is an e_mux
  assign cpu_instruction_master_read_data_valid_epcs_epcs_control_port = cpu_instruction_master_granted_epcs_epcs_control_port & cpu_instruction_master_read & ~epcs_epcs_control_port_waits_for_read;

  //allow new arb cycle for epcs/epcs_control_port, which is an e_assign
  assign epcs_epcs_control_port_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock;

  //cpu/instruction_master assignment into master qualified-requests vector for epcs/epcs_control_port, which is an e_assign
  assign epcs_epcs_control_port_master_qreq_vector[0] = cpu_instruction_master_qualified_request_epcs_epcs_control_port;

  //cpu/instruction_master grant epcs/epcs_control_port, which is an e_assign
  assign cpu_instruction_master_granted_epcs_epcs_control_port = epcs_epcs_control_port_grant_vector[0];

  //cpu/instruction_master saved-grant epcs/epcs_control_port, which is an e_assign
  assign cpu_instruction_master_saved_grant_epcs_epcs_control_port = epcs_epcs_control_port_arb_winner[0] && cpu_instruction_master_requests_epcs_epcs_control_port;

  //cpu/data_master assignment into master qualified-requests vector for epcs/epcs_control_port, which is an e_assign
  assign epcs_epcs_control_port_master_qreq_vector[1] = cpu_data_master_qualified_request_epcs_epcs_control_port;

  //cpu/data_master grant epcs/epcs_control_port, which is an e_assign
  assign cpu_data_master_granted_epcs_epcs_control_port = epcs_epcs_control_port_grant_vector[1];

  //cpu/data_master saved-grant epcs/epcs_control_port, which is an e_assign
  assign cpu_data_master_saved_grant_epcs_epcs_control_port = epcs_epcs_control_port_arb_winner[1] && cpu_data_master_requests_epcs_epcs_control_port;

  //epcs/epcs_control_port chosen-master double-vector, which is an e_assign
  assign epcs_epcs_control_port_chosen_master_double_vector = {epcs_epcs_control_port_master_qreq_vector, epcs_epcs_control_port_master_qreq_vector} & ({~epcs_epcs_control_port_master_qreq_vector, ~epcs_epcs_control_port_master_qreq_vector} + epcs_epcs_control_port_arb_addend);

  //stable onehot encoding of arb winner
  assign epcs_epcs_control_port_arb_winner = (epcs_epcs_control_port_allow_new_arb_cycle & | epcs_epcs_control_port_grant_vector) ? epcs_epcs_control_port_grant_vector : epcs_epcs_control_port_saved_chosen_master_vector;

  //saved epcs_epcs_control_port_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          epcs_epcs_control_port_saved_chosen_master_vector <= 0;
      else if (epcs_epcs_control_port_allow_new_arb_cycle)
          epcs_epcs_control_port_saved_chosen_master_vector <= |epcs_epcs_control_port_grant_vector ? epcs_epcs_control_port_grant_vector : epcs_epcs_control_port_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign epcs_epcs_control_port_grant_vector = {(epcs_epcs_control_port_chosen_master_double_vector[1] | epcs_epcs_control_port_chosen_master_double_vector[3]),
    (epcs_epcs_control_port_chosen_master_double_vector[0] | epcs_epcs_control_port_chosen_master_double_vector[2])};

  //epcs/epcs_control_port chosen master rotated left, which is an e_assign
  assign epcs_epcs_control_port_chosen_master_rot_left = (epcs_epcs_control_port_arb_winner << 1) ? (epcs_epcs_control_port_arb_winner << 1) : 1;

  //epcs/epcs_control_port's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          epcs_epcs_control_port_arb_addend <= 1;
      else if (|epcs_epcs_control_port_grant_vector)
          epcs_epcs_control_port_arb_addend <= epcs_epcs_control_port_end_xfer? epcs_epcs_control_port_chosen_master_rot_left : epcs_epcs_control_port_grant_vector;
    end


  //epcs_epcs_control_port_reset_n assignment, which is an e_assign
  assign epcs_epcs_control_port_reset_n = reset_n;

  assign epcs_epcs_control_port_chipselect = cpu_data_master_granted_epcs_epcs_control_port | cpu_instruction_master_granted_epcs_epcs_control_port;
  //epcs_epcs_control_port_firsttransfer first transaction, which is an e_assign
  assign epcs_epcs_control_port_firsttransfer = epcs_epcs_control_port_begins_xfer ? epcs_epcs_control_port_unreg_firsttransfer : epcs_epcs_control_port_reg_firsttransfer;

  //epcs_epcs_control_port_unreg_firsttransfer first transaction, which is an e_assign
  assign epcs_epcs_control_port_unreg_firsttransfer = ~(epcs_epcs_control_port_slavearbiterlockenable & epcs_epcs_control_port_any_continuerequest);

  //epcs_epcs_control_port_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          epcs_epcs_control_port_reg_firsttransfer <= 1'b1;
      else if (epcs_epcs_control_port_begins_xfer)
          epcs_epcs_control_port_reg_firsttransfer <= epcs_epcs_control_port_unreg_firsttransfer;
    end


  //epcs_epcs_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign epcs_epcs_control_port_beginbursttransfer_internal = epcs_epcs_control_port_begins_xfer;

  //epcs_epcs_control_port_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign epcs_epcs_control_port_arbitration_holdoff_internal = epcs_epcs_control_port_begins_xfer & epcs_epcs_control_port_firsttransfer;

  //~epcs_epcs_control_port_read_n assignment, which is an e_mux
  assign epcs_epcs_control_port_read_n = ~((cpu_data_master_granted_epcs_epcs_control_port & cpu_data_master_read) | (cpu_instruction_master_granted_epcs_epcs_control_port & cpu_instruction_master_read));

  //~epcs_epcs_control_port_write_n assignment, which is an e_mux
  assign epcs_epcs_control_port_write_n = ~(cpu_data_master_granted_epcs_epcs_control_port & cpu_data_master_write);

  assign shifted_address_to_epcs_epcs_control_port_from_cpu_data_master = cpu_data_master_address_to_slave;
  //epcs_epcs_control_port_address mux, which is an e_mux
  assign epcs_epcs_control_port_address = (cpu_data_master_granted_epcs_epcs_control_port)? (shifted_address_to_epcs_epcs_control_port_from_cpu_data_master >> 2) :
    (shifted_address_to_epcs_epcs_control_port_from_cpu_instruction_master >> 2);

  assign shifted_address_to_epcs_epcs_control_port_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  //d1_epcs_epcs_control_port_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_epcs_epcs_control_port_end_xfer <= 1;
      else 
        d1_epcs_epcs_control_port_end_xfer <= epcs_epcs_control_port_end_xfer;
    end


  //epcs_epcs_control_port_waits_for_read in a cycle, which is an e_mux
  assign epcs_epcs_control_port_waits_for_read = epcs_epcs_control_port_in_a_read_cycle & epcs_epcs_control_port_begins_xfer;

  //epcs_epcs_control_port_in_a_read_cycle assignment, which is an e_assign
  assign epcs_epcs_control_port_in_a_read_cycle = (cpu_data_master_granted_epcs_epcs_control_port & cpu_data_master_read) | (cpu_instruction_master_granted_epcs_epcs_control_port & cpu_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = epcs_epcs_control_port_in_a_read_cycle;

  //epcs_epcs_control_port_waits_for_write in a cycle, which is an e_mux
  assign epcs_epcs_control_port_waits_for_write = epcs_epcs_control_port_in_a_write_cycle & epcs_epcs_control_port_begins_xfer;

  //epcs_epcs_control_port_in_a_write_cycle assignment, which is an e_assign
  assign epcs_epcs_control_port_in_a_write_cycle = cpu_data_master_granted_epcs_epcs_control_port & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = epcs_epcs_control_port_in_a_write_cycle;

  assign wait_for_epcs_epcs_control_port_counter = 0;
  //assign epcs_epcs_control_port_irq_from_sa = epcs_epcs_control_port_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign epcs_epcs_control_port_irq_from_sa = epcs_epcs_control_port_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //epcs/epcs_control_port enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_epcs_epcs_control_port + cpu_instruction_master_granted_epcs_epcs_control_port > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_epcs_epcs_control_port + cpu_instruction_master_saved_grant_epcs_epcs_control_port > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_avalon_jtag_slave_arbitrator (
                                                // inputs:
                                                 clk,
                                                 cpu_data_master_address_to_slave,
                                                 cpu_data_master_read,
                                                 cpu_data_master_waitrequest,
                                                 cpu_data_master_write,
                                                 cpu_data_master_writedata,
                                                 jtag_uart_avalon_jtag_slave_dataavailable,
                                                 jtag_uart_avalon_jtag_slave_irq,
                                                 jtag_uart_avalon_jtag_slave_readdata,
                                                 jtag_uart_avalon_jtag_slave_readyfordata,
                                                 jtag_uart_avalon_jtag_slave_waitrequest,
                                                 reset_n,

                                                // outputs:
                                                 cpu_data_master_granted_jtag_uart_avalon_jtag_slave,
                                                 cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave,
                                                 cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave,
                                                 cpu_data_master_requests_jtag_uart_avalon_jtag_slave,
                                                 d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                                 jtag_uart_avalon_jtag_slave_address,
                                                 jtag_uart_avalon_jtag_slave_chipselect,
                                                 jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
                                                 jtag_uart_avalon_jtag_slave_irq_from_sa,
                                                 jtag_uart_avalon_jtag_slave_read_n,
                                                 jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_reset_n,
                                                 jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                                 jtag_uart_avalon_jtag_slave_write_n,
                                                 jtag_uart_avalon_jtag_slave_writedata
                                              )
;

  output           cpu_data_master_granted_jtag_uart_avalon_jtag_slave;
  output           cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave;
  output           cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave;
  output           cpu_data_master_requests_jtag_uart_avalon_jtag_slave;
  output           d1_jtag_uart_avalon_jtag_slave_end_xfer;
  output           jtag_uart_avalon_jtag_slave_address;
  output           jtag_uart_avalon_jtag_slave_chipselect;
  output           jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_avalon_jtag_slave_reset_n;
  output           jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_read;
  input            cpu_data_master_waitrequest;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            jtag_uart_avalon_jtag_slave_dataavailable;
  input            jtag_uart_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  input            jtag_uart_avalon_jtag_slave_readyfordata;
  input            jtag_uart_avalon_jtag_slave_waitrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_requests_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_saved_grant_jtag_uart_avalon_jtag_slave;
  reg              d1_jtag_uart_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_allgrants;
  wire             jtag_uart_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_avalon_jtag_slave_arb_counter_enable;
  reg     [  1: 0] jtag_uart_avalon_jtag_slave_arb_share_counter;
  wire    [  1: 0] jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
  wire    [  1: 0] jtag_uart_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  reg              jtag_uart_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire    [ 26: 0] shifted_address_to_jtag_uart_avalon_jtag_slave_from_cpu_data_master;
  wire             wait_for_jtag_uart_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~jtag_uart_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave));
  //assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata;

  assign cpu_data_master_requests_jtag_uart_avalon_jtag_slave = ({cpu_data_master_address_to_slave[26 : 3] , 3'b0} == 27'h1898) & (cpu_data_master_read | cpu_data_master_write);
  //assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest;

  //jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_arb_share_set_values = 1;

  //jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_non_bursting_master_requests = cpu_data_master_requests_jtag_uart_avalon_jtag_slave;

  //jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant = 0;

  //jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_avalon_jtag_slave_firsttransfer ? (jtag_uart_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_avalon_jtag_slave_arb_share_counter ? (jtag_uart_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_allgrants = |jtag_uart_avalon_jtag_slave_grant_vector;

  //jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_end_xfer = ~(jtag_uart_avalon_jtag_slave_waits_for_read | jtag_uart_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave = jtag_uart_avalon_jtag_slave_end_xfer & (~jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & jtag_uart_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //cpu/data_master jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = jtag_uart_avalon_jtag_slave_slavearbiterlockenable & cpu_data_master_continuerequest;

  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;

  //cpu/data_master jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave = cpu_data_master_requests_jtag_uart_avalon_jtag_slave & ~((cpu_data_master_read & (~cpu_data_master_waitrequest)) | ((~cpu_data_master_waitrequest) & cpu_data_master_write));
  //jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_jtag_uart_avalon_jtag_slave = cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave;

  //cpu/data_master saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  assign cpu_data_master_saved_grant_jtag_uart_avalon_jtag_slave = cpu_data_master_requests_jtag_uart_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_avalon_jtag_slave_chipselect = cpu_data_master_granted_jtag_uart_avalon_jtag_slave;
  //jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_firsttransfer = jtag_uart_avalon_jtag_slave_begins_xfer ? jtag_uart_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_avalon_jtag_slave_begins_xfer)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_read_n = ~(cpu_data_master_granted_jtag_uart_avalon_jtag_slave & cpu_data_master_read);

  //~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_write_n = ~(cpu_data_master_granted_jtag_uart_avalon_jtag_slave & cpu_data_master_write);

  assign shifted_address_to_jtag_uart_avalon_jtag_slave_from_cpu_data_master = cpu_data_master_address_to_slave;
  //jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_address = shifted_address_to_jtag_uart_avalon_jtag_slave_from_cpu_data_master >> 2;

  //d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_avalon_jtag_slave_end_xfer <= 1;
      else 
        d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_read = jtag_uart_avalon_jtag_slave_in_a_read_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_read_cycle = cpu_data_master_granted_jtag_uart_avalon_jtag_slave & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_write = jtag_uart_avalon_jtag_slave_in_a_write_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_write_cycle = cpu_data_master_granted_jtag_uart_avalon_jtag_slave & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_sdram_s1_module (
                                                         // inputs:
                                                          clear_fifo,
                                                          clk,
                                                          data_in,
                                                          read,
                                                          reset_n,
                                                          sync_reset,
                                                          write,

                                                         // outputs:
                                                          data_out,
                                                          empty,
                                                          fifo_contains_ones_n,
                                                          full
                                                       )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  wire             full_6;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_5;
  assign empty = !full_0;
  assign full_6 = 0;
  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    0;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_sdram_s1_module (
                                                                // inputs:
                                                                 clear_fifo,
                                                                 clk,
                                                                 data_in,
                                                                 read,
                                                                 reset_n,
                                                                 sync_reset,
                                                                 write,

                                                                // outputs:
                                                                 data_out,
                                                                 empty,
                                                                 fifo_contains_ones_n,
                                                                 full
                                                              )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  wire             full_6;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_5;
  assign empty = !full_0;
  assign full_6 = 0;
  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    0;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sdram_s1_arbitrator (
                             // inputs:
                              clk,
                              cpu_data_master_address_to_slave,
                              cpu_data_master_byteenable,
                              cpu_data_master_dbs_address,
                              cpu_data_master_dbs_write_16,
                              cpu_data_master_no_byte_enables_and_last_term,
                              cpu_data_master_read,
                              cpu_data_master_waitrequest,
                              cpu_data_master_write,
                              cpu_instruction_master_address_to_slave,
                              cpu_instruction_master_dbs_address,
                              cpu_instruction_master_latency_counter,
                              cpu_instruction_master_read,
                              reset_n,
                              sdram_s1_readdata,
                              sdram_s1_readdatavalid,
                              sdram_s1_waitrequest,

                             // outputs:
                              cpu_data_master_byteenable_sdram_s1,
                              cpu_data_master_granted_sdram_s1,
                              cpu_data_master_qualified_request_sdram_s1,
                              cpu_data_master_read_data_valid_sdram_s1,
                              cpu_data_master_read_data_valid_sdram_s1_shift_register,
                              cpu_data_master_requests_sdram_s1,
                              cpu_instruction_master_granted_sdram_s1,
                              cpu_instruction_master_qualified_request_sdram_s1,
                              cpu_instruction_master_read_data_valid_sdram_s1,
                              cpu_instruction_master_read_data_valid_sdram_s1_shift_register,
                              cpu_instruction_master_requests_sdram_s1,
                              d1_sdram_s1_end_xfer,
                              sdram_s1_address,
                              sdram_s1_byteenable_n,
                              sdram_s1_chipselect,
                              sdram_s1_read_n,
                              sdram_s1_readdata_from_sa,
                              sdram_s1_reset_n,
                              sdram_s1_waitrequest_from_sa,
                              sdram_s1_write_n,
                              sdram_s1_writedata
                           )
;

  output  [  1: 0] cpu_data_master_byteenable_sdram_s1;
  output           cpu_data_master_granted_sdram_s1;
  output           cpu_data_master_qualified_request_sdram_s1;
  output           cpu_data_master_read_data_valid_sdram_s1;
  output           cpu_data_master_read_data_valid_sdram_s1_shift_register;
  output           cpu_data_master_requests_sdram_s1;
  output           cpu_instruction_master_granted_sdram_s1;
  output           cpu_instruction_master_qualified_request_sdram_s1;
  output           cpu_instruction_master_read_data_valid_sdram_s1;
  output           cpu_instruction_master_read_data_valid_sdram_s1_shift_register;
  output           cpu_instruction_master_requests_sdram_s1;
  output           d1_sdram_s1_end_xfer;
  output  [ 23: 0] sdram_s1_address;
  output  [  1: 0] sdram_s1_byteenable_n;
  output           sdram_s1_chipselect;
  output           sdram_s1_read_n;
  output  [ 15: 0] sdram_s1_readdata_from_sa;
  output           sdram_s1_reset_n;
  output           sdram_s1_waitrequest_from_sa;
  output           sdram_s1_write_n;
  output  [ 15: 0] sdram_s1_writedata;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input   [  1: 0] cpu_data_master_dbs_address;
  input   [ 15: 0] cpu_data_master_dbs_write_16;
  input            cpu_data_master_no_byte_enables_and_last_term;
  input            cpu_data_master_read;
  input            cpu_data_master_waitrequest;
  input            cpu_data_master_write;
  input   [ 26: 0] cpu_instruction_master_address_to_slave;
  input   [  1: 0] cpu_instruction_master_dbs_address;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            reset_n;
  input   [ 15: 0] sdram_s1_readdata;
  input            sdram_s1_readdatavalid;
  input            sdram_s1_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire    [  1: 0] cpu_data_master_byteenable_sdram_s1;
  wire    [  1: 0] cpu_data_master_byteenable_sdram_s1_segment_0;
  wire    [  1: 0] cpu_data_master_byteenable_sdram_s1_segment_1;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_sdram_s1;
  wire             cpu_data_master_qualified_request_sdram_s1;
  wire             cpu_data_master_rdv_fifo_empty_sdram_s1;
  wire             cpu_data_master_rdv_fifo_output_from_sdram_s1;
  wire             cpu_data_master_read_data_valid_sdram_s1;
  wire             cpu_data_master_read_data_valid_sdram_s1_shift_register;
  wire             cpu_data_master_requests_sdram_s1;
  wire             cpu_data_master_saved_grant_sdram_s1;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_sdram_s1;
  wire             cpu_instruction_master_qualified_request_sdram_s1;
  wire             cpu_instruction_master_rdv_fifo_empty_sdram_s1;
  wire             cpu_instruction_master_rdv_fifo_output_from_sdram_s1;
  wire             cpu_instruction_master_read_data_valid_sdram_s1;
  wire             cpu_instruction_master_read_data_valid_sdram_s1_shift_register;
  wire             cpu_instruction_master_requests_sdram_s1;
  wire             cpu_instruction_master_saved_grant_sdram_s1;
  reg              d1_reasons_to_wait;
  reg              d1_sdram_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sdram_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_sdram_s1;
  reg              last_cycle_cpu_instruction_master_granted_slave_sdram_s1;
  wire    [ 23: 0] sdram_s1_address;
  wire             sdram_s1_allgrants;
  wire             sdram_s1_allow_new_arb_cycle;
  wire             sdram_s1_any_bursting_master_saved_grant;
  wire             sdram_s1_any_continuerequest;
  reg     [  1: 0] sdram_s1_arb_addend;
  wire             sdram_s1_arb_counter_enable;
  reg     [  1: 0] sdram_s1_arb_share_counter;
  wire    [  1: 0] sdram_s1_arb_share_counter_next_value;
  wire    [  1: 0] sdram_s1_arb_share_set_values;
  wire    [  1: 0] sdram_s1_arb_winner;
  wire             sdram_s1_arbitration_holdoff_internal;
  wire             sdram_s1_beginbursttransfer_internal;
  wire             sdram_s1_begins_xfer;
  wire    [  1: 0] sdram_s1_byteenable_n;
  wire             sdram_s1_chipselect;
  wire    [  3: 0] sdram_s1_chosen_master_double_vector;
  wire    [  1: 0] sdram_s1_chosen_master_rot_left;
  wire             sdram_s1_end_xfer;
  wire             sdram_s1_firsttransfer;
  wire    [  1: 0] sdram_s1_grant_vector;
  wire             sdram_s1_in_a_read_cycle;
  wire             sdram_s1_in_a_write_cycle;
  wire    [  1: 0] sdram_s1_master_qreq_vector;
  wire             sdram_s1_move_on_to_next_transaction;
  wire             sdram_s1_non_bursting_master_requests;
  wire             sdram_s1_read_n;
  wire    [ 15: 0] sdram_s1_readdata_from_sa;
  wire             sdram_s1_readdatavalid_from_sa;
  reg              sdram_s1_reg_firsttransfer;
  wire             sdram_s1_reset_n;
  reg     [  1: 0] sdram_s1_saved_chosen_master_vector;
  reg              sdram_s1_slavearbiterlockenable;
  wire             sdram_s1_slavearbiterlockenable2;
  wire             sdram_s1_unreg_firsttransfer;
  wire             sdram_s1_waitrequest_from_sa;
  wire             sdram_s1_waits_for_read;
  wire             sdram_s1_waits_for_write;
  wire             sdram_s1_write_n;
  wire    [ 15: 0] sdram_s1_writedata;
  wire    [ 26: 0] shifted_address_to_sdram_s1_from_cpu_data_master;
  wire    [ 26: 0] shifted_address_to_sdram_s1_from_cpu_instruction_master;
  wire             wait_for_sdram_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sdram_s1_end_xfer;
    end


  assign sdram_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_sdram_s1 | cpu_instruction_master_qualified_request_sdram_s1));
  //assign sdram_s1_readdatavalid_from_sa = sdram_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sdram_s1_readdatavalid_from_sa = sdram_s1_readdatavalid;

  //assign sdram_s1_readdata_from_sa = sdram_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sdram_s1_readdata_from_sa = sdram_s1_readdata;

  assign cpu_data_master_requests_sdram_s1 = ({cpu_data_master_address_to_slave[26 : 25] , 25'b0} == 27'h4000000) & (cpu_data_master_read | cpu_data_master_write);
  //assign sdram_s1_waitrequest_from_sa = sdram_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sdram_s1_waitrequest_from_sa = sdram_s1_waitrequest;

  //sdram_s1_arb_share_counter set values, which is an e_mux
  assign sdram_s1_arb_share_set_values = (cpu_data_master_granted_sdram_s1)? 2 :
    (cpu_instruction_master_granted_sdram_s1)? 2 :
    (cpu_data_master_granted_sdram_s1)? 2 :
    (cpu_instruction_master_granted_sdram_s1)? 2 :
    1;

  //sdram_s1_non_bursting_master_requests mux, which is an e_mux
  assign sdram_s1_non_bursting_master_requests = cpu_data_master_requests_sdram_s1 |
    cpu_instruction_master_requests_sdram_s1 |
    cpu_data_master_requests_sdram_s1 |
    cpu_instruction_master_requests_sdram_s1;

  //sdram_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign sdram_s1_any_bursting_master_saved_grant = 0;

  //sdram_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign sdram_s1_arb_share_counter_next_value = sdram_s1_firsttransfer ? (sdram_s1_arb_share_set_values - 1) : |sdram_s1_arb_share_counter ? (sdram_s1_arb_share_counter - 1) : 0;

  //sdram_s1_allgrants all slave grants, which is an e_mux
  assign sdram_s1_allgrants = (|sdram_s1_grant_vector) |
    (|sdram_s1_grant_vector) |
    (|sdram_s1_grant_vector) |
    (|sdram_s1_grant_vector);

  //sdram_s1_end_xfer assignment, which is an e_assign
  assign sdram_s1_end_xfer = ~(sdram_s1_waits_for_read | sdram_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_sdram_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sdram_s1 = sdram_s1_end_xfer & (~sdram_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sdram_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign sdram_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_sdram_s1 & sdram_s1_allgrants) | (end_xfer_arb_share_counter_term_sdram_s1 & ~sdram_s1_non_bursting_master_requests);

  //sdram_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_s1_arb_share_counter <= 0;
      else if (sdram_s1_arb_counter_enable)
          sdram_s1_arb_share_counter <= sdram_s1_arb_share_counter_next_value;
    end


  //sdram_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_s1_slavearbiterlockenable <= 0;
      else if ((|sdram_s1_master_qreq_vector & end_xfer_arb_share_counter_term_sdram_s1) | (end_xfer_arb_share_counter_term_sdram_s1 & ~sdram_s1_non_bursting_master_requests))
          sdram_s1_slavearbiterlockenable <= |sdram_s1_arb_share_counter_next_value;
    end


  //cpu/data_master sdram/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = sdram_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //sdram_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sdram_s1_slavearbiterlockenable2 = |sdram_s1_arb_share_counter_next_value;

  //cpu/data_master sdram/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = sdram_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master sdram/s1 arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = sdram_s1_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master sdram/s1 arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = sdram_s1_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted sdram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_sdram_s1 <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_sdram_s1 <= cpu_instruction_master_saved_grant_sdram_s1 ? 1 : (sdram_s1_arbitration_holdoff_internal | ~cpu_instruction_master_requests_sdram_s1) ? 0 : last_cycle_cpu_instruction_master_granted_slave_sdram_s1;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = last_cycle_cpu_instruction_master_granted_slave_sdram_s1 & cpu_instruction_master_requests_sdram_s1;

  //sdram_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign sdram_s1_any_continuerequest = cpu_instruction_master_continuerequest |
    cpu_data_master_continuerequest;

  assign cpu_data_master_qualified_request_sdram_s1 = cpu_data_master_requests_sdram_s1 & ~((cpu_data_master_read & (~cpu_data_master_waitrequest | (|cpu_data_master_read_data_valid_sdram_s1_shift_register))) | ((~cpu_data_master_waitrequest | cpu_data_master_no_byte_enables_and_last_term | !cpu_data_master_byteenable_sdram_s1) & cpu_data_master_write) | cpu_instruction_master_arbiterlock);
  //unique name for sdram_s1_move_on_to_next_transaction, which is an e_assign
  assign sdram_s1_move_on_to_next_transaction = sdram_s1_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_sdram_s1_module rdv_fifo_for_cpu_data_master_to_sdram_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_sdram_s1),
      .data_out             (cpu_data_master_rdv_fifo_output_from_sdram_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_sdram_s1),
      .full                 (),
      .read                 (sdram_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_s1_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_sdram_s1_shift_register = ~cpu_data_master_rdv_fifo_empty_sdram_s1;
  //local readdatavalid cpu_data_master_read_data_valid_sdram_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_sdram_s1 = (sdram_s1_readdatavalid_from_sa & cpu_data_master_rdv_fifo_output_from_sdram_s1) & ~ cpu_data_master_rdv_fifo_empty_sdram_s1;

  //sdram_s1_writedata mux, which is an e_mux
  assign sdram_s1_writedata = cpu_data_master_dbs_write_16;

  assign cpu_instruction_master_requests_sdram_s1 = (({cpu_instruction_master_address_to_slave[26 : 25] , 25'b0} == 27'h4000000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted sdram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_sdram_s1 <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_sdram_s1 <= cpu_data_master_saved_grant_sdram_s1 ? 1 : (sdram_s1_arbitration_holdoff_internal | ~cpu_data_master_requests_sdram_s1) ? 0 : last_cycle_cpu_data_master_granted_slave_sdram_s1;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = last_cycle_cpu_data_master_granted_slave_sdram_s1 & cpu_data_master_requests_sdram_s1;

  assign cpu_instruction_master_qualified_request_sdram_s1 = cpu_instruction_master_requests_sdram_s1 & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter))) | cpu_data_master_arbiterlock);
  //rdv_fifo_for_cpu_instruction_master_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_sdram_s1_module rdv_fifo_for_cpu_instruction_master_to_sdram_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_sdram_s1),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_sdram_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_sdram_s1),
      .full                 (),
      .read                 (sdram_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_s1_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_sdram_s1_shift_register = ~cpu_instruction_master_rdv_fifo_empty_sdram_s1;
  //local readdatavalid cpu_instruction_master_read_data_valid_sdram_s1, which is an e_mux
  assign cpu_instruction_master_read_data_valid_sdram_s1 = (sdram_s1_readdatavalid_from_sa & cpu_instruction_master_rdv_fifo_output_from_sdram_s1) & ~ cpu_instruction_master_rdv_fifo_empty_sdram_s1;

  //allow new arb cycle for sdram/s1, which is an e_assign
  assign sdram_s1_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock;

  //cpu/instruction_master assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  assign sdram_s1_master_qreq_vector[0] = cpu_instruction_master_qualified_request_sdram_s1;

  //cpu/instruction_master grant sdram/s1, which is an e_assign
  assign cpu_instruction_master_granted_sdram_s1 = sdram_s1_grant_vector[0];

  //cpu/instruction_master saved-grant sdram/s1, which is an e_assign
  assign cpu_instruction_master_saved_grant_sdram_s1 = sdram_s1_arb_winner[0] && cpu_instruction_master_requests_sdram_s1;

  //cpu/data_master assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  assign sdram_s1_master_qreq_vector[1] = cpu_data_master_qualified_request_sdram_s1;

  //cpu/data_master grant sdram/s1, which is an e_assign
  assign cpu_data_master_granted_sdram_s1 = sdram_s1_grant_vector[1];

  //cpu/data_master saved-grant sdram/s1, which is an e_assign
  assign cpu_data_master_saved_grant_sdram_s1 = sdram_s1_arb_winner[1] && cpu_data_master_requests_sdram_s1;

  //sdram/s1 chosen-master double-vector, which is an e_assign
  assign sdram_s1_chosen_master_double_vector = {sdram_s1_master_qreq_vector, sdram_s1_master_qreq_vector} & ({~sdram_s1_master_qreq_vector, ~sdram_s1_master_qreq_vector} + sdram_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign sdram_s1_arb_winner = (sdram_s1_allow_new_arb_cycle & | sdram_s1_grant_vector) ? sdram_s1_grant_vector : sdram_s1_saved_chosen_master_vector;

  //saved sdram_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_s1_saved_chosen_master_vector <= 0;
      else if (sdram_s1_allow_new_arb_cycle)
          sdram_s1_saved_chosen_master_vector <= |sdram_s1_grant_vector ? sdram_s1_grant_vector : sdram_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign sdram_s1_grant_vector = {(sdram_s1_chosen_master_double_vector[1] | sdram_s1_chosen_master_double_vector[3]),
    (sdram_s1_chosen_master_double_vector[0] | sdram_s1_chosen_master_double_vector[2])};

  //sdram/s1 chosen master rotated left, which is an e_assign
  assign sdram_s1_chosen_master_rot_left = (sdram_s1_arb_winner << 1) ? (sdram_s1_arb_winner << 1) : 1;

  //sdram/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_s1_arb_addend <= 1;
      else if (|sdram_s1_grant_vector)
          sdram_s1_arb_addend <= sdram_s1_end_xfer? sdram_s1_chosen_master_rot_left : sdram_s1_grant_vector;
    end


  //sdram_s1_reset_n assignment, which is an e_assign
  assign sdram_s1_reset_n = reset_n;

  assign sdram_s1_chipselect = cpu_data_master_granted_sdram_s1 | cpu_instruction_master_granted_sdram_s1;
  //sdram_s1_firsttransfer first transaction, which is an e_assign
  assign sdram_s1_firsttransfer = sdram_s1_begins_xfer ? sdram_s1_unreg_firsttransfer : sdram_s1_reg_firsttransfer;

  //sdram_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign sdram_s1_unreg_firsttransfer = ~(sdram_s1_slavearbiterlockenable & sdram_s1_any_continuerequest);

  //sdram_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_s1_reg_firsttransfer <= 1'b1;
      else if (sdram_s1_begins_xfer)
          sdram_s1_reg_firsttransfer <= sdram_s1_unreg_firsttransfer;
    end


  //sdram_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sdram_s1_beginbursttransfer_internal = sdram_s1_begins_xfer;

  //sdram_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign sdram_s1_arbitration_holdoff_internal = sdram_s1_begins_xfer & sdram_s1_firsttransfer;

  //~sdram_s1_read_n assignment, which is an e_mux
  assign sdram_s1_read_n = ~((cpu_data_master_granted_sdram_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_sdram_s1 & cpu_instruction_master_read));

  //~sdram_s1_write_n assignment, which is an e_mux
  assign sdram_s1_write_n = ~(cpu_data_master_granted_sdram_s1 & cpu_data_master_write);

  assign shifted_address_to_sdram_s1_from_cpu_data_master = {cpu_data_master_address_to_slave >> 2,
    cpu_data_master_dbs_address[1],
    {1 {1'b0}}};

  //sdram_s1_address mux, which is an e_mux
  assign sdram_s1_address = (cpu_data_master_granted_sdram_s1)? (shifted_address_to_sdram_s1_from_cpu_data_master >> 1) :
    (shifted_address_to_sdram_s1_from_cpu_instruction_master >> 1);

  assign shifted_address_to_sdram_s1_from_cpu_instruction_master = {cpu_instruction_master_address_to_slave >> 2,
    cpu_instruction_master_dbs_address[1],
    {1 {1'b0}}};

  //d1_sdram_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sdram_s1_end_xfer <= 1;
      else 
        d1_sdram_s1_end_xfer <= sdram_s1_end_xfer;
    end


  //sdram_s1_waits_for_read in a cycle, which is an e_mux
  assign sdram_s1_waits_for_read = sdram_s1_in_a_read_cycle & sdram_s1_waitrequest_from_sa;

  //sdram_s1_in_a_read_cycle assignment, which is an e_assign
  assign sdram_s1_in_a_read_cycle = (cpu_data_master_granted_sdram_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_sdram_s1 & cpu_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sdram_s1_in_a_read_cycle;

  //sdram_s1_waits_for_write in a cycle, which is an e_mux
  assign sdram_s1_waits_for_write = sdram_s1_in_a_write_cycle & sdram_s1_waitrequest_from_sa;

  //sdram_s1_in_a_write_cycle assignment, which is an e_assign
  assign sdram_s1_in_a_write_cycle = cpu_data_master_granted_sdram_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sdram_s1_in_a_write_cycle;

  assign wait_for_sdram_s1_counter = 0;
  //~sdram_s1_byteenable_n byte enable port mux, which is an e_mux
  assign sdram_s1_byteenable_n = ~((cpu_data_master_granted_sdram_s1)? cpu_data_master_byteenable_sdram_s1 :
    -1);

  assign {cpu_data_master_byteenable_sdram_s1_segment_1,
cpu_data_master_byteenable_sdram_s1_segment_0} = cpu_data_master_byteenable;
  assign cpu_data_master_byteenable_sdram_s1 = ((cpu_data_master_dbs_address[1] == 0))? cpu_data_master_byteenable_sdram_s1_segment_0 :
    cpu_data_master_byteenable_sdram_s1_segment_1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sdram/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_sdram_s1 + cpu_instruction_master_granted_sdram_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_sdram_s1 + cpu_instruction_master_saved_grant_sdram_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sysid_control_slave_arbitrator (
                                        // inputs:
                                         clk,
                                         cpu_data_master_address_to_slave,
                                         cpu_data_master_read,
                                         cpu_data_master_write,
                                         reset_n,
                                         sysid_control_slave_readdata,

                                        // outputs:
                                         cpu_data_master_granted_sysid_control_slave,
                                         cpu_data_master_qualified_request_sysid_control_slave,
                                         cpu_data_master_read_data_valid_sysid_control_slave,
                                         cpu_data_master_requests_sysid_control_slave,
                                         d1_sysid_control_slave_end_xfer,
                                         sysid_control_slave_address,
                                         sysid_control_slave_readdata_from_sa,
                                         sysid_control_slave_reset_n
                                      )
;

  output           cpu_data_master_granted_sysid_control_slave;
  output           cpu_data_master_qualified_request_sysid_control_slave;
  output           cpu_data_master_read_data_valid_sysid_control_slave;
  output           cpu_data_master_requests_sysid_control_slave;
  output           d1_sysid_control_slave_end_xfer;
  output           sysid_control_slave_address;
  output  [ 31: 0] sysid_control_slave_readdata_from_sa;
  output           sysid_control_slave_reset_n;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_read;
  input            cpu_data_master_write;
  input            reset_n;
  input   [ 31: 0] sysid_control_slave_readdata;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_sysid_control_slave;
  wire             cpu_data_master_qualified_request_sysid_control_slave;
  wire             cpu_data_master_read_data_valid_sysid_control_slave;
  wire             cpu_data_master_requests_sysid_control_slave;
  wire             cpu_data_master_saved_grant_sysid_control_slave;
  reg              d1_reasons_to_wait;
  reg              d1_sysid_control_slave_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sysid_control_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 26: 0] shifted_address_to_sysid_control_slave_from_cpu_data_master;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_allgrants;
  wire             sysid_control_slave_allow_new_arb_cycle;
  wire             sysid_control_slave_any_bursting_master_saved_grant;
  wire             sysid_control_slave_any_continuerequest;
  wire             sysid_control_slave_arb_counter_enable;
  reg     [  1: 0] sysid_control_slave_arb_share_counter;
  wire    [  1: 0] sysid_control_slave_arb_share_counter_next_value;
  wire    [  1: 0] sysid_control_slave_arb_share_set_values;
  wire             sysid_control_slave_beginbursttransfer_internal;
  wire             sysid_control_slave_begins_xfer;
  wire             sysid_control_slave_end_xfer;
  wire             sysid_control_slave_firsttransfer;
  wire             sysid_control_slave_grant_vector;
  wire             sysid_control_slave_in_a_read_cycle;
  wire             sysid_control_slave_in_a_write_cycle;
  wire             sysid_control_slave_master_qreq_vector;
  wire             sysid_control_slave_non_bursting_master_requests;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  reg              sysid_control_slave_reg_firsttransfer;
  wire             sysid_control_slave_reset_n;
  reg              sysid_control_slave_slavearbiterlockenable;
  wire             sysid_control_slave_slavearbiterlockenable2;
  wire             sysid_control_slave_unreg_firsttransfer;
  wire             sysid_control_slave_waits_for_read;
  wire             sysid_control_slave_waits_for_write;
  wire             wait_for_sysid_control_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sysid_control_slave_end_xfer;
    end


  assign sysid_control_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_sysid_control_slave));
  //assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata;

  assign cpu_data_master_requests_sysid_control_slave = (({cpu_data_master_address_to_slave[26 : 3] , 3'b0} == 27'h1890) & (cpu_data_master_read | cpu_data_master_write)) & cpu_data_master_read;
  //sysid_control_slave_arb_share_counter set values, which is an e_mux
  assign sysid_control_slave_arb_share_set_values = 1;

  //sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  assign sysid_control_slave_non_bursting_master_requests = cpu_data_master_requests_sysid_control_slave;

  //sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign sysid_control_slave_any_bursting_master_saved_grant = 0;

  //sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign sysid_control_slave_arb_share_counter_next_value = sysid_control_slave_firsttransfer ? (sysid_control_slave_arb_share_set_values - 1) : |sysid_control_slave_arb_share_counter ? (sysid_control_slave_arb_share_counter - 1) : 0;

  //sysid_control_slave_allgrants all slave grants, which is an e_mux
  assign sysid_control_slave_allgrants = |sysid_control_slave_grant_vector;

  //sysid_control_slave_end_xfer assignment, which is an e_assign
  assign sysid_control_slave_end_xfer = ~(sysid_control_slave_waits_for_read | sysid_control_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sysid_control_slave = sysid_control_slave_end_xfer & (~sysid_control_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign sysid_control_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_sysid_control_slave & sysid_control_slave_allgrants) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests);

  //sysid_control_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_arb_share_counter <= 0;
      else if (sysid_control_slave_arb_counter_enable)
          sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
    end


  //sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_slavearbiterlockenable <= 0;
      else if ((|sysid_control_slave_master_qreq_vector & end_xfer_arb_share_counter_term_sysid_control_slave) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests))
          sysid_control_slave_slavearbiterlockenable <= |sysid_control_slave_arb_share_counter_next_value;
    end


  //cpu/data_master sysid/control_slave arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = sysid_control_slave_slavearbiterlockenable & cpu_data_master_continuerequest;

  //sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sysid_control_slave_slavearbiterlockenable2 = |sysid_control_slave_arb_share_counter_next_value;

  //cpu/data_master sysid/control_slave arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = sysid_control_slave_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sysid_control_slave_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_sysid_control_slave = cpu_data_master_requests_sysid_control_slave;
  //master is always granted when requested
  assign cpu_data_master_granted_sysid_control_slave = cpu_data_master_qualified_request_sysid_control_slave;

  //cpu/data_master saved-grant sysid/control_slave, which is an e_assign
  assign cpu_data_master_saved_grant_sysid_control_slave = cpu_data_master_requests_sysid_control_slave;

  //allow new arb cycle for sysid/control_slave, which is an e_assign
  assign sysid_control_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sysid_control_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sysid_control_slave_master_qreq_vector = 1;

  //sysid_control_slave_reset_n assignment, which is an e_assign
  assign sysid_control_slave_reset_n = reset_n;

  //sysid_control_slave_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_firsttransfer = sysid_control_slave_begins_xfer ? sysid_control_slave_unreg_firsttransfer : sysid_control_slave_reg_firsttransfer;

  //sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_unreg_firsttransfer = ~(sysid_control_slave_slavearbiterlockenable & sysid_control_slave_any_continuerequest);

  //sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_reg_firsttransfer <= 1'b1;
      else if (sysid_control_slave_begins_xfer)
          sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
    end


  //sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sysid_control_slave_beginbursttransfer_internal = sysid_control_slave_begins_xfer;

  assign shifted_address_to_sysid_control_slave_from_cpu_data_master = cpu_data_master_address_to_slave;
  //sysid_control_slave_address mux, which is an e_mux
  assign sysid_control_slave_address = shifted_address_to_sysid_control_slave_from_cpu_data_master >> 2;

  //d1_sysid_control_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sysid_control_slave_end_xfer <= 1;
      else 
        d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end


  //sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_read = sysid_control_slave_in_a_read_cycle & sysid_control_slave_begins_xfer;

  //sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_read_cycle = cpu_data_master_granted_sysid_control_slave & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sysid_control_slave_in_a_read_cycle;

  //sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_write = sysid_control_slave_in_a_write_cycle & 0;

  //sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_write_cycle = cpu_data_master_granted_sysid_control_slave & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sysid_control_slave_in_a_write_cycle;

  assign wait_for_sysid_control_slave_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sysid/control_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module kernel_reset_clk_domain_synch_module (
                                              // inputs:
                                               clk,
                                               data_in,
                                               reset_n,

                                              // outputs:
                                               data_out
                                            )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module kernel (
                // 1) global signals:
                 clk,
                 reset_n,

                // the_PIO_LCD_B
                 out_port_from_the_PIO_LCD_B,

                // the_PIO_LCD_CLK
                 out_port_from_the_PIO_LCD_CLK,

                // the_PIO_LCD_CTRL
                 out_port_from_the_PIO_LCD_CTRL,

                // the_PIO_LCD_G
                 out_port_from_the_PIO_LCD_G,

                // the_PIO_LCD_PWM
                 out_port_from_the_PIO_LCD_PWM,

                // the_PIO_LCD_R
                 out_port_from_the_PIO_LCD_R,

                // the_PIO_LED
                 out_port_from_the_PIO_LED,

                // the_RS232
                 rxd_to_the_RS232,
                 txd_from_the_RS232,

                // the_epcs
                 data0_to_the_epcs,
                 dclk_from_the_epcs,
                 sce_from_the_epcs,
                 sdo_from_the_epcs,

                // the_sdram
                 zs_addr_from_the_sdram,
                 zs_ba_from_the_sdram,
                 zs_cas_n_from_the_sdram,
                 zs_cke_from_the_sdram,
                 zs_cs_n_from_the_sdram,
                 zs_dq_to_and_from_the_sdram,
                 zs_dqm_from_the_sdram,
                 zs_ras_n_from_the_sdram,
                 zs_we_n_from_the_sdram
              )
;

  output           dclk_from_the_epcs;
  output  [  5: 0] out_port_from_the_PIO_LCD_B;
  output           out_port_from_the_PIO_LCD_CLK;
  output  [  7: 0] out_port_from_the_PIO_LCD_CTRL;
  output  [  5: 0] out_port_from_the_PIO_LCD_G;
  output           out_port_from_the_PIO_LCD_PWM;
  output  [  5: 0] out_port_from_the_PIO_LCD_R;
  output  [  3: 0] out_port_from_the_PIO_LED;
  output           sce_from_the_epcs;
  output           sdo_from_the_epcs;
  output           txd_from_the_RS232;
  output  [ 12: 0] zs_addr_from_the_sdram;
  output  [  1: 0] zs_ba_from_the_sdram;
  output           zs_cas_n_from_the_sdram;
  output           zs_cke_from_the_sdram;
  output           zs_cs_n_from_the_sdram;
  inout   [ 15: 0] zs_dq_to_and_from_the_sdram;
  output  [  1: 0] zs_dqm_from_the_sdram;
  output           zs_ras_n_from_the_sdram;
  output           zs_we_n_from_the_sdram;
  input            clk;
  input            data0_to_the_epcs;
  input            reset_n;
  input            rxd_to_the_RS232;

  wire    [  1: 0] PIO_LCD_B_s1_address;
  wire             PIO_LCD_B_s1_chipselect;
  wire    [ 31: 0] PIO_LCD_B_s1_readdata;
  wire    [ 31: 0] PIO_LCD_B_s1_readdata_from_sa;
  wire             PIO_LCD_B_s1_reset_n;
  wire             PIO_LCD_B_s1_write_n;
  wire    [ 31: 0] PIO_LCD_B_s1_writedata;
  wire    [  1: 0] PIO_LCD_CLK_s1_address;
  wire             PIO_LCD_CLK_s1_chipselect;
  wire    [ 31: 0] PIO_LCD_CLK_s1_readdata;
  wire    [ 31: 0] PIO_LCD_CLK_s1_readdata_from_sa;
  wire             PIO_LCD_CLK_s1_reset_n;
  wire             PIO_LCD_CLK_s1_write_n;
  wire    [ 31: 0] PIO_LCD_CLK_s1_writedata;
  wire    [  1: 0] PIO_LCD_CTRL_s1_address;
  wire             PIO_LCD_CTRL_s1_chipselect;
  wire    [ 31: 0] PIO_LCD_CTRL_s1_readdata;
  wire    [ 31: 0] PIO_LCD_CTRL_s1_readdata_from_sa;
  wire             PIO_LCD_CTRL_s1_reset_n;
  wire             PIO_LCD_CTRL_s1_write_n;
  wire    [ 31: 0] PIO_LCD_CTRL_s1_writedata;
  wire    [  1: 0] PIO_LCD_G_s1_address;
  wire             PIO_LCD_G_s1_chipselect;
  wire    [ 31: 0] PIO_LCD_G_s1_readdata;
  wire    [ 31: 0] PIO_LCD_G_s1_readdata_from_sa;
  wire             PIO_LCD_G_s1_reset_n;
  wire             PIO_LCD_G_s1_write_n;
  wire    [ 31: 0] PIO_LCD_G_s1_writedata;
  wire    [  1: 0] PIO_LCD_PWM_s1_address;
  wire             PIO_LCD_PWM_s1_chipselect;
  wire    [ 31: 0] PIO_LCD_PWM_s1_readdata;
  wire    [ 31: 0] PIO_LCD_PWM_s1_readdata_from_sa;
  wire             PIO_LCD_PWM_s1_reset_n;
  wire             PIO_LCD_PWM_s1_write_n;
  wire    [ 31: 0] PIO_LCD_PWM_s1_writedata;
  wire    [  1: 0] PIO_LCD_R_s1_address;
  wire             PIO_LCD_R_s1_chipselect;
  wire    [ 31: 0] PIO_LCD_R_s1_readdata;
  wire    [ 31: 0] PIO_LCD_R_s1_readdata_from_sa;
  wire             PIO_LCD_R_s1_reset_n;
  wire             PIO_LCD_R_s1_write_n;
  wire    [ 31: 0] PIO_LCD_R_s1_writedata;
  wire    [  1: 0] PIO_LED_s1_address;
  wire             PIO_LED_s1_chipselect;
  wire    [ 31: 0] PIO_LED_s1_readdata;
  wire    [ 31: 0] PIO_LED_s1_readdata_from_sa;
  wire             PIO_LED_s1_reset_n;
  wire             PIO_LED_s1_write_n;
  wire    [ 31: 0] PIO_LED_s1_writedata;
  wire    [  2: 0] RS232_s1_address;
  wire             RS232_s1_begintransfer;
  wire             RS232_s1_chipselect;
  wire             RS232_s1_dataavailable;
  wire             RS232_s1_dataavailable_from_sa;
  wire             RS232_s1_irq;
  wire             RS232_s1_irq_from_sa;
  wire             RS232_s1_read_n;
  wire    [ 15: 0] RS232_s1_readdata;
  wire    [ 15: 0] RS232_s1_readdata_from_sa;
  wire             RS232_s1_readyfordata;
  wire             RS232_s1_readyfordata_from_sa;
  wire             RS232_s1_reset_n;
  wire             RS232_s1_write_n;
  wire    [ 15: 0] RS232_s1_writedata;
  wire             clk_reset_n;
  wire    [ 26: 0] cpu_data_master_address;
  wire    [ 26: 0] cpu_data_master_address_to_slave;
  wire    [  3: 0] cpu_data_master_byteenable;
  wire    [  1: 0] cpu_data_master_byteenable_sdram_s1;
  wire    [  1: 0] cpu_data_master_dbs_address;
  wire    [ 15: 0] cpu_data_master_dbs_write_16;
  wire             cpu_data_master_debugaccess;
  wire             cpu_data_master_granted_PIO_LCD_B_s1;
  wire             cpu_data_master_granted_PIO_LCD_CLK_s1;
  wire             cpu_data_master_granted_PIO_LCD_CTRL_s1;
  wire             cpu_data_master_granted_PIO_LCD_G_s1;
  wire             cpu_data_master_granted_PIO_LCD_PWM_s1;
  wire             cpu_data_master_granted_PIO_LCD_R_s1;
  wire             cpu_data_master_granted_PIO_LED_s1;
  wire             cpu_data_master_granted_RS232_s1;
  wire             cpu_data_master_granted_cpu_jtag_debug_module;
  wire             cpu_data_master_granted_epcs_epcs_control_port;
  wire             cpu_data_master_granted_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_granted_sdram_s1;
  wire             cpu_data_master_granted_sysid_control_slave;
  wire    [ 31: 0] cpu_data_master_irq;
  wire             cpu_data_master_no_byte_enables_and_last_term;
  wire             cpu_data_master_qualified_request_PIO_LCD_B_s1;
  wire             cpu_data_master_qualified_request_PIO_LCD_CLK_s1;
  wire             cpu_data_master_qualified_request_PIO_LCD_CTRL_s1;
  wire             cpu_data_master_qualified_request_PIO_LCD_G_s1;
  wire             cpu_data_master_qualified_request_PIO_LCD_PWM_s1;
  wire             cpu_data_master_qualified_request_PIO_LCD_R_s1;
  wire             cpu_data_master_qualified_request_PIO_LED_s1;
  wire             cpu_data_master_qualified_request_RS232_s1;
  wire             cpu_data_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_data_master_qualified_request_epcs_epcs_control_port;
  wire             cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_qualified_request_sdram_s1;
  wire             cpu_data_master_qualified_request_sysid_control_slave;
  wire             cpu_data_master_read;
  wire             cpu_data_master_read_data_valid_PIO_LCD_B_s1;
  wire             cpu_data_master_read_data_valid_PIO_LCD_CLK_s1;
  wire             cpu_data_master_read_data_valid_PIO_LCD_CTRL_s1;
  wire             cpu_data_master_read_data_valid_PIO_LCD_G_s1;
  wire             cpu_data_master_read_data_valid_PIO_LCD_PWM_s1;
  wire             cpu_data_master_read_data_valid_PIO_LCD_R_s1;
  wire             cpu_data_master_read_data_valid_PIO_LED_s1;
  wire             cpu_data_master_read_data_valid_RS232_s1;
  wire             cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_data_master_read_data_valid_epcs_epcs_control_port;
  wire             cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_read_data_valid_sdram_s1;
  wire             cpu_data_master_read_data_valid_sdram_s1_shift_register;
  wire             cpu_data_master_read_data_valid_sysid_control_slave;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_requests_PIO_LCD_B_s1;
  wire             cpu_data_master_requests_PIO_LCD_CLK_s1;
  wire             cpu_data_master_requests_PIO_LCD_CTRL_s1;
  wire             cpu_data_master_requests_PIO_LCD_G_s1;
  wire             cpu_data_master_requests_PIO_LCD_PWM_s1;
  wire             cpu_data_master_requests_PIO_LCD_R_s1;
  wire             cpu_data_master_requests_PIO_LED_s1;
  wire             cpu_data_master_requests_RS232_s1;
  wire             cpu_data_master_requests_cpu_jtag_debug_module;
  wire             cpu_data_master_requests_epcs_epcs_control_port;
  wire             cpu_data_master_requests_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_requests_sdram_s1;
  wire             cpu_data_master_requests_sysid_control_slave;
  wire             cpu_data_master_waitrequest;
  wire             cpu_data_master_write;
  wire    [ 31: 0] cpu_data_master_writedata;
  wire    [ 26: 0] cpu_instruction_master_address;
  wire    [ 26: 0] cpu_instruction_master_address_to_slave;
  wire    [  1: 0] cpu_instruction_master_dbs_address;
  wire             cpu_instruction_master_granted_cpu_jtag_debug_module;
  wire             cpu_instruction_master_granted_epcs_epcs_control_port;
  wire             cpu_instruction_master_granted_sdram_s1;
  wire             cpu_instruction_master_latency_counter;
  wire             cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_instruction_master_qualified_request_epcs_epcs_control_port;
  wire             cpu_instruction_master_qualified_request_sdram_s1;
  wire             cpu_instruction_master_read;
  wire             cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_instruction_master_read_data_valid_epcs_epcs_control_port;
  wire             cpu_instruction_master_read_data_valid_sdram_s1;
  wire             cpu_instruction_master_read_data_valid_sdram_s1_shift_register;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_requests_cpu_jtag_debug_module;
  wire             cpu_instruction_master_requests_epcs_epcs_control_port;
  wire             cpu_instruction_master_requests_sdram_s1;
  wire             cpu_instruction_master_waitrequest;
  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire             cpu_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  wire             d1_PIO_LCD_B_s1_end_xfer;
  wire             d1_PIO_LCD_CLK_s1_end_xfer;
  wire             d1_PIO_LCD_CTRL_s1_end_xfer;
  wire             d1_PIO_LCD_G_s1_end_xfer;
  wire             d1_PIO_LCD_PWM_s1_end_xfer;
  wire             d1_PIO_LCD_R_s1_end_xfer;
  wire             d1_PIO_LED_s1_end_xfer;
  wire             d1_RS232_s1_end_xfer;
  wire             d1_cpu_jtag_debug_module_end_xfer;
  wire             d1_epcs_epcs_control_port_end_xfer;
  wire             d1_jtag_uart_avalon_jtag_slave_end_xfer;
  wire             d1_sdram_s1_end_xfer;
  wire             d1_sysid_control_slave_end_xfer;
  wire             dclk_from_the_epcs;
  wire    [  8: 0] epcs_epcs_control_port_address;
  wire             epcs_epcs_control_port_chipselect;
  wire             epcs_epcs_control_port_dataavailable;
  wire             epcs_epcs_control_port_dataavailable_from_sa;
  wire             epcs_epcs_control_port_endofpacket;
  wire             epcs_epcs_control_port_endofpacket_from_sa;
  wire             epcs_epcs_control_port_irq;
  wire             epcs_epcs_control_port_irq_from_sa;
  wire             epcs_epcs_control_port_read_n;
  wire    [ 31: 0] epcs_epcs_control_port_readdata;
  wire    [ 31: 0] epcs_epcs_control_port_readdata_from_sa;
  wire             epcs_epcs_control_port_readyfordata;
  wire             epcs_epcs_control_port_readyfordata_from_sa;
  wire             epcs_epcs_control_port_reset_n;
  wire             epcs_epcs_control_port_write_n;
  wire    [ 31: 0] epcs_epcs_control_port_writedata;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_irq;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  wire             jtag_uart_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire    [  5: 0] out_port_from_the_PIO_LCD_B;
  wire             out_port_from_the_PIO_LCD_CLK;
  wire    [  7: 0] out_port_from_the_PIO_LCD_CTRL;
  wire    [  5: 0] out_port_from_the_PIO_LCD_G;
  wire             out_port_from_the_PIO_LCD_PWM;
  wire    [  5: 0] out_port_from_the_PIO_LCD_R;
  wire    [  3: 0] out_port_from_the_PIO_LED;
  wire             reset_n_sources;
  wire             sce_from_the_epcs;
  wire             sdo_from_the_epcs;
  wire    [ 23: 0] sdram_s1_address;
  wire    [  1: 0] sdram_s1_byteenable_n;
  wire             sdram_s1_chipselect;
  wire             sdram_s1_read_n;
  wire    [ 15: 0] sdram_s1_readdata;
  wire    [ 15: 0] sdram_s1_readdata_from_sa;
  wire             sdram_s1_readdatavalid;
  wire             sdram_s1_reset_n;
  wire             sdram_s1_waitrequest;
  wire             sdram_s1_waitrequest_from_sa;
  wire             sdram_s1_write_n;
  wire    [ 15: 0] sdram_s1_writedata;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_clock;
  wire    [ 31: 0] sysid_control_slave_readdata;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  wire             sysid_control_slave_reset_n;
  wire             txd_from_the_RS232;
  wire    [ 12: 0] zs_addr_from_the_sdram;
  wire    [  1: 0] zs_ba_from_the_sdram;
  wire             zs_cas_n_from_the_sdram;
  wire             zs_cke_from_the_sdram;
  wire             zs_cs_n_from_the_sdram;
  wire    [ 15: 0] zs_dq_to_and_from_the_sdram;
  wire    [  1: 0] zs_dqm_from_the_sdram;
  wire             zs_ras_n_from_the_sdram;
  wire             zs_we_n_from_the_sdram;
  PIO_LCD_B_s1_arbitrator the_PIO_LCD_B_s1
    (
      .PIO_LCD_B_s1_address                           (PIO_LCD_B_s1_address),
      .PIO_LCD_B_s1_chipselect                        (PIO_LCD_B_s1_chipselect),
      .PIO_LCD_B_s1_readdata                          (PIO_LCD_B_s1_readdata),
      .PIO_LCD_B_s1_readdata_from_sa                  (PIO_LCD_B_s1_readdata_from_sa),
      .PIO_LCD_B_s1_reset_n                           (PIO_LCD_B_s1_reset_n),
      .PIO_LCD_B_s1_write_n                           (PIO_LCD_B_s1_write_n),
      .PIO_LCD_B_s1_writedata                         (PIO_LCD_B_s1_writedata),
      .clk                                            (clk),
      .cpu_data_master_address_to_slave               (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_PIO_LCD_B_s1           (cpu_data_master_granted_PIO_LCD_B_s1),
      .cpu_data_master_qualified_request_PIO_LCD_B_s1 (cpu_data_master_qualified_request_PIO_LCD_B_s1),
      .cpu_data_master_read                           (cpu_data_master_read),
      .cpu_data_master_read_data_valid_PIO_LCD_B_s1   (cpu_data_master_read_data_valid_PIO_LCD_B_s1),
      .cpu_data_master_requests_PIO_LCD_B_s1          (cpu_data_master_requests_PIO_LCD_B_s1),
      .cpu_data_master_waitrequest                    (cpu_data_master_waitrequest),
      .cpu_data_master_write                          (cpu_data_master_write),
      .cpu_data_master_writedata                      (cpu_data_master_writedata),
      .d1_PIO_LCD_B_s1_end_xfer                       (d1_PIO_LCD_B_s1_end_xfer),
      .reset_n                                        (clk_reset_n)
    );

  PIO_LCD_B the_PIO_LCD_B
    (
      .address    (PIO_LCD_B_s1_address),
      .chipselect (PIO_LCD_B_s1_chipselect),
      .clk        (clk),
      .out_port   (out_port_from_the_PIO_LCD_B),
      .readdata   (PIO_LCD_B_s1_readdata),
      .reset_n    (PIO_LCD_B_s1_reset_n),
      .write_n    (PIO_LCD_B_s1_write_n),
      .writedata  (PIO_LCD_B_s1_writedata)
    );

  PIO_LCD_CLK_s1_arbitrator the_PIO_LCD_CLK_s1
    (
      .PIO_LCD_CLK_s1_address                           (PIO_LCD_CLK_s1_address),
      .PIO_LCD_CLK_s1_chipselect                        (PIO_LCD_CLK_s1_chipselect),
      .PIO_LCD_CLK_s1_readdata                          (PIO_LCD_CLK_s1_readdata),
      .PIO_LCD_CLK_s1_readdata_from_sa                  (PIO_LCD_CLK_s1_readdata_from_sa),
      .PIO_LCD_CLK_s1_reset_n                           (PIO_LCD_CLK_s1_reset_n),
      .PIO_LCD_CLK_s1_write_n                           (PIO_LCD_CLK_s1_write_n),
      .PIO_LCD_CLK_s1_writedata                         (PIO_LCD_CLK_s1_writedata),
      .clk                                              (clk),
      .cpu_data_master_address_to_slave                 (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_PIO_LCD_CLK_s1           (cpu_data_master_granted_PIO_LCD_CLK_s1),
      .cpu_data_master_qualified_request_PIO_LCD_CLK_s1 (cpu_data_master_qualified_request_PIO_LCD_CLK_s1),
      .cpu_data_master_read                             (cpu_data_master_read),
      .cpu_data_master_read_data_valid_PIO_LCD_CLK_s1   (cpu_data_master_read_data_valid_PIO_LCD_CLK_s1),
      .cpu_data_master_requests_PIO_LCD_CLK_s1          (cpu_data_master_requests_PIO_LCD_CLK_s1),
      .cpu_data_master_waitrequest                      (cpu_data_master_waitrequest),
      .cpu_data_master_write                            (cpu_data_master_write),
      .cpu_data_master_writedata                        (cpu_data_master_writedata),
      .d1_PIO_LCD_CLK_s1_end_xfer                       (d1_PIO_LCD_CLK_s1_end_xfer),
      .reset_n                                          (clk_reset_n)
    );

  PIO_LCD_CLK the_PIO_LCD_CLK
    (
      .address    (PIO_LCD_CLK_s1_address),
      .chipselect (PIO_LCD_CLK_s1_chipselect),
      .clk        (clk),
      .out_port   (out_port_from_the_PIO_LCD_CLK),
      .readdata   (PIO_LCD_CLK_s1_readdata),
      .reset_n    (PIO_LCD_CLK_s1_reset_n),
      .write_n    (PIO_LCD_CLK_s1_write_n),
      .writedata  (PIO_LCD_CLK_s1_writedata)
    );

  PIO_LCD_CTRL_s1_arbitrator the_PIO_LCD_CTRL_s1
    (
      .PIO_LCD_CTRL_s1_address                           (PIO_LCD_CTRL_s1_address),
      .PIO_LCD_CTRL_s1_chipselect                        (PIO_LCD_CTRL_s1_chipselect),
      .PIO_LCD_CTRL_s1_readdata                          (PIO_LCD_CTRL_s1_readdata),
      .PIO_LCD_CTRL_s1_readdata_from_sa                  (PIO_LCD_CTRL_s1_readdata_from_sa),
      .PIO_LCD_CTRL_s1_reset_n                           (PIO_LCD_CTRL_s1_reset_n),
      .PIO_LCD_CTRL_s1_write_n                           (PIO_LCD_CTRL_s1_write_n),
      .PIO_LCD_CTRL_s1_writedata                         (PIO_LCD_CTRL_s1_writedata),
      .clk                                               (clk),
      .cpu_data_master_address_to_slave                  (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_PIO_LCD_CTRL_s1           (cpu_data_master_granted_PIO_LCD_CTRL_s1),
      .cpu_data_master_qualified_request_PIO_LCD_CTRL_s1 (cpu_data_master_qualified_request_PIO_LCD_CTRL_s1),
      .cpu_data_master_read                              (cpu_data_master_read),
      .cpu_data_master_read_data_valid_PIO_LCD_CTRL_s1   (cpu_data_master_read_data_valid_PIO_LCD_CTRL_s1),
      .cpu_data_master_requests_PIO_LCD_CTRL_s1          (cpu_data_master_requests_PIO_LCD_CTRL_s1),
      .cpu_data_master_waitrequest                       (cpu_data_master_waitrequest),
      .cpu_data_master_write                             (cpu_data_master_write),
      .cpu_data_master_writedata                         (cpu_data_master_writedata),
      .d1_PIO_LCD_CTRL_s1_end_xfer                       (d1_PIO_LCD_CTRL_s1_end_xfer),
      .reset_n                                           (clk_reset_n)
    );

  PIO_LCD_CTRL the_PIO_LCD_CTRL
    (
      .address    (PIO_LCD_CTRL_s1_address),
      .chipselect (PIO_LCD_CTRL_s1_chipselect),
      .clk        (clk),
      .out_port   (out_port_from_the_PIO_LCD_CTRL),
      .readdata   (PIO_LCD_CTRL_s1_readdata),
      .reset_n    (PIO_LCD_CTRL_s1_reset_n),
      .write_n    (PIO_LCD_CTRL_s1_write_n),
      .writedata  (PIO_LCD_CTRL_s1_writedata)
    );

  PIO_LCD_G_s1_arbitrator the_PIO_LCD_G_s1
    (
      .PIO_LCD_G_s1_address                           (PIO_LCD_G_s1_address),
      .PIO_LCD_G_s1_chipselect                        (PIO_LCD_G_s1_chipselect),
      .PIO_LCD_G_s1_readdata                          (PIO_LCD_G_s1_readdata),
      .PIO_LCD_G_s1_readdata_from_sa                  (PIO_LCD_G_s1_readdata_from_sa),
      .PIO_LCD_G_s1_reset_n                           (PIO_LCD_G_s1_reset_n),
      .PIO_LCD_G_s1_write_n                           (PIO_LCD_G_s1_write_n),
      .PIO_LCD_G_s1_writedata                         (PIO_LCD_G_s1_writedata),
      .clk                                            (clk),
      .cpu_data_master_address_to_slave               (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_PIO_LCD_G_s1           (cpu_data_master_granted_PIO_LCD_G_s1),
      .cpu_data_master_qualified_request_PIO_LCD_G_s1 (cpu_data_master_qualified_request_PIO_LCD_G_s1),
      .cpu_data_master_read                           (cpu_data_master_read),
      .cpu_data_master_read_data_valid_PIO_LCD_G_s1   (cpu_data_master_read_data_valid_PIO_LCD_G_s1),
      .cpu_data_master_requests_PIO_LCD_G_s1          (cpu_data_master_requests_PIO_LCD_G_s1),
      .cpu_data_master_waitrequest                    (cpu_data_master_waitrequest),
      .cpu_data_master_write                          (cpu_data_master_write),
      .cpu_data_master_writedata                      (cpu_data_master_writedata),
      .d1_PIO_LCD_G_s1_end_xfer                       (d1_PIO_LCD_G_s1_end_xfer),
      .reset_n                                        (clk_reset_n)
    );

  PIO_LCD_G the_PIO_LCD_G
    (
      .address    (PIO_LCD_G_s1_address),
      .chipselect (PIO_LCD_G_s1_chipselect),
      .clk        (clk),
      .out_port   (out_port_from_the_PIO_LCD_G),
      .readdata   (PIO_LCD_G_s1_readdata),
      .reset_n    (PIO_LCD_G_s1_reset_n),
      .write_n    (PIO_LCD_G_s1_write_n),
      .writedata  (PIO_LCD_G_s1_writedata)
    );

  PIO_LCD_PWM_s1_arbitrator the_PIO_LCD_PWM_s1
    (
      .PIO_LCD_PWM_s1_address                           (PIO_LCD_PWM_s1_address),
      .PIO_LCD_PWM_s1_chipselect                        (PIO_LCD_PWM_s1_chipselect),
      .PIO_LCD_PWM_s1_readdata                          (PIO_LCD_PWM_s1_readdata),
      .PIO_LCD_PWM_s1_readdata_from_sa                  (PIO_LCD_PWM_s1_readdata_from_sa),
      .PIO_LCD_PWM_s1_reset_n                           (PIO_LCD_PWM_s1_reset_n),
      .PIO_LCD_PWM_s1_write_n                           (PIO_LCD_PWM_s1_write_n),
      .PIO_LCD_PWM_s1_writedata                         (PIO_LCD_PWM_s1_writedata),
      .clk                                              (clk),
      .cpu_data_master_address_to_slave                 (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_PIO_LCD_PWM_s1           (cpu_data_master_granted_PIO_LCD_PWM_s1),
      .cpu_data_master_qualified_request_PIO_LCD_PWM_s1 (cpu_data_master_qualified_request_PIO_LCD_PWM_s1),
      .cpu_data_master_read                             (cpu_data_master_read),
      .cpu_data_master_read_data_valid_PIO_LCD_PWM_s1   (cpu_data_master_read_data_valid_PIO_LCD_PWM_s1),
      .cpu_data_master_requests_PIO_LCD_PWM_s1          (cpu_data_master_requests_PIO_LCD_PWM_s1),
      .cpu_data_master_waitrequest                      (cpu_data_master_waitrequest),
      .cpu_data_master_write                            (cpu_data_master_write),
      .cpu_data_master_writedata                        (cpu_data_master_writedata),
      .d1_PIO_LCD_PWM_s1_end_xfer                       (d1_PIO_LCD_PWM_s1_end_xfer),
      .reset_n                                          (clk_reset_n)
    );

  PIO_LCD_PWM the_PIO_LCD_PWM
    (
      .address    (PIO_LCD_PWM_s1_address),
      .chipselect (PIO_LCD_PWM_s1_chipselect),
      .clk        (clk),
      .out_port   (out_port_from_the_PIO_LCD_PWM),
      .readdata   (PIO_LCD_PWM_s1_readdata),
      .reset_n    (PIO_LCD_PWM_s1_reset_n),
      .write_n    (PIO_LCD_PWM_s1_write_n),
      .writedata  (PIO_LCD_PWM_s1_writedata)
    );

  PIO_LCD_R_s1_arbitrator the_PIO_LCD_R_s1
    (
      .PIO_LCD_R_s1_address                           (PIO_LCD_R_s1_address),
      .PIO_LCD_R_s1_chipselect                        (PIO_LCD_R_s1_chipselect),
      .PIO_LCD_R_s1_readdata                          (PIO_LCD_R_s1_readdata),
      .PIO_LCD_R_s1_readdata_from_sa                  (PIO_LCD_R_s1_readdata_from_sa),
      .PIO_LCD_R_s1_reset_n                           (PIO_LCD_R_s1_reset_n),
      .PIO_LCD_R_s1_write_n                           (PIO_LCD_R_s1_write_n),
      .PIO_LCD_R_s1_writedata                         (PIO_LCD_R_s1_writedata),
      .clk                                            (clk),
      .cpu_data_master_address_to_slave               (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_PIO_LCD_R_s1           (cpu_data_master_granted_PIO_LCD_R_s1),
      .cpu_data_master_qualified_request_PIO_LCD_R_s1 (cpu_data_master_qualified_request_PIO_LCD_R_s1),
      .cpu_data_master_read                           (cpu_data_master_read),
      .cpu_data_master_read_data_valid_PIO_LCD_R_s1   (cpu_data_master_read_data_valid_PIO_LCD_R_s1),
      .cpu_data_master_requests_PIO_LCD_R_s1          (cpu_data_master_requests_PIO_LCD_R_s1),
      .cpu_data_master_waitrequest                    (cpu_data_master_waitrequest),
      .cpu_data_master_write                          (cpu_data_master_write),
      .cpu_data_master_writedata                      (cpu_data_master_writedata),
      .d1_PIO_LCD_R_s1_end_xfer                       (d1_PIO_LCD_R_s1_end_xfer),
      .reset_n                                        (clk_reset_n)
    );

  PIO_LCD_R the_PIO_LCD_R
    (
      .address    (PIO_LCD_R_s1_address),
      .chipselect (PIO_LCD_R_s1_chipselect),
      .clk        (clk),
      .out_port   (out_port_from_the_PIO_LCD_R),
      .readdata   (PIO_LCD_R_s1_readdata),
      .reset_n    (PIO_LCD_R_s1_reset_n),
      .write_n    (PIO_LCD_R_s1_write_n),
      .writedata  (PIO_LCD_R_s1_writedata)
    );

  PIO_LED_s1_arbitrator the_PIO_LED_s1
    (
      .PIO_LED_s1_address                           (PIO_LED_s1_address),
      .PIO_LED_s1_chipselect                        (PIO_LED_s1_chipselect),
      .PIO_LED_s1_readdata                          (PIO_LED_s1_readdata),
      .PIO_LED_s1_readdata_from_sa                  (PIO_LED_s1_readdata_from_sa),
      .PIO_LED_s1_reset_n                           (PIO_LED_s1_reset_n),
      .PIO_LED_s1_write_n                           (PIO_LED_s1_write_n),
      .PIO_LED_s1_writedata                         (PIO_LED_s1_writedata),
      .clk                                          (clk),
      .cpu_data_master_address_to_slave             (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_PIO_LED_s1           (cpu_data_master_granted_PIO_LED_s1),
      .cpu_data_master_qualified_request_PIO_LED_s1 (cpu_data_master_qualified_request_PIO_LED_s1),
      .cpu_data_master_read                         (cpu_data_master_read),
      .cpu_data_master_read_data_valid_PIO_LED_s1   (cpu_data_master_read_data_valid_PIO_LED_s1),
      .cpu_data_master_requests_PIO_LED_s1          (cpu_data_master_requests_PIO_LED_s1),
      .cpu_data_master_waitrequest                  (cpu_data_master_waitrequest),
      .cpu_data_master_write                        (cpu_data_master_write),
      .cpu_data_master_writedata                    (cpu_data_master_writedata),
      .d1_PIO_LED_s1_end_xfer                       (d1_PIO_LED_s1_end_xfer),
      .reset_n                                      (clk_reset_n)
    );

  PIO_LED the_PIO_LED
    (
      .address    (PIO_LED_s1_address),
      .chipselect (PIO_LED_s1_chipselect),
      .clk        (clk),
      .out_port   (out_port_from_the_PIO_LED),
      .readdata   (PIO_LED_s1_readdata),
      .reset_n    (PIO_LED_s1_reset_n),
      .write_n    (PIO_LED_s1_write_n),
      .writedata  (PIO_LED_s1_writedata)
    );

  RS232_s1_arbitrator the_RS232_s1
    (
      .RS232_s1_address                           (RS232_s1_address),
      .RS232_s1_begintransfer                     (RS232_s1_begintransfer),
      .RS232_s1_chipselect                        (RS232_s1_chipselect),
      .RS232_s1_dataavailable                     (RS232_s1_dataavailable),
      .RS232_s1_dataavailable_from_sa             (RS232_s1_dataavailable_from_sa),
      .RS232_s1_irq                               (RS232_s1_irq),
      .RS232_s1_irq_from_sa                       (RS232_s1_irq_from_sa),
      .RS232_s1_read_n                            (RS232_s1_read_n),
      .RS232_s1_readdata                          (RS232_s1_readdata),
      .RS232_s1_readdata_from_sa                  (RS232_s1_readdata_from_sa),
      .RS232_s1_readyfordata                      (RS232_s1_readyfordata),
      .RS232_s1_readyfordata_from_sa              (RS232_s1_readyfordata_from_sa),
      .RS232_s1_reset_n                           (RS232_s1_reset_n),
      .RS232_s1_write_n                           (RS232_s1_write_n),
      .RS232_s1_writedata                         (RS232_s1_writedata),
      .clk                                        (clk),
      .cpu_data_master_address_to_slave           (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_RS232_s1           (cpu_data_master_granted_RS232_s1),
      .cpu_data_master_qualified_request_RS232_s1 (cpu_data_master_qualified_request_RS232_s1),
      .cpu_data_master_read                       (cpu_data_master_read),
      .cpu_data_master_read_data_valid_RS232_s1   (cpu_data_master_read_data_valid_RS232_s1),
      .cpu_data_master_requests_RS232_s1          (cpu_data_master_requests_RS232_s1),
      .cpu_data_master_write                      (cpu_data_master_write),
      .cpu_data_master_writedata                  (cpu_data_master_writedata),
      .d1_RS232_s1_end_xfer                       (d1_RS232_s1_end_xfer),
      .reset_n                                    (clk_reset_n)
    );

  RS232 the_RS232
    (
      .address       (RS232_s1_address),
      .begintransfer (RS232_s1_begintransfer),
      .chipselect    (RS232_s1_chipselect),
      .clk           (clk),
      .dataavailable (RS232_s1_dataavailable),
      .irq           (RS232_s1_irq),
      .read_n        (RS232_s1_read_n),
      .readdata      (RS232_s1_readdata),
      .readyfordata  (RS232_s1_readyfordata),
      .reset_n       (RS232_s1_reset_n),
      .rxd           (rxd_to_the_RS232),
      .txd           (txd_from_the_RS232),
      .write_n       (RS232_s1_write_n),
      .writedata     (RS232_s1_writedata)
    );

  cpu_jtag_debug_module_arbitrator the_cpu_jtag_debug_module
    (
      .clk                                                            (clk),
      .cpu_data_master_address_to_slave                               (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                     (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                    (cpu_data_master_debugaccess),
      .cpu_data_master_granted_cpu_jtag_debug_module                  (cpu_data_master_granted_cpu_jtag_debug_module),
      .cpu_data_master_qualified_request_cpu_jtag_debug_module        (cpu_data_master_qualified_request_cpu_jtag_debug_module),
      .cpu_data_master_read                                           (cpu_data_master_read),
      .cpu_data_master_read_data_valid_cpu_jtag_debug_module          (cpu_data_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_data_master_requests_cpu_jtag_debug_module                 (cpu_data_master_requests_cpu_jtag_debug_module),
      .cpu_data_master_waitrequest                                    (cpu_data_master_waitrequest),
      .cpu_data_master_write                                          (cpu_data_master_write),
      .cpu_data_master_writedata                                      (cpu_data_master_writedata),
      .cpu_instruction_master_address_to_slave                        (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_cpu_jtag_debug_module           (cpu_instruction_master_granted_cpu_jtag_debug_module),
      .cpu_instruction_master_latency_counter                         (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_cpu_jtag_debug_module (cpu_instruction_master_qualified_request_cpu_jtag_debug_module),
      .cpu_instruction_master_read                                    (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_cpu_jtag_debug_module   (cpu_instruction_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_instruction_master_read_data_valid_sdram_s1_shift_register (cpu_instruction_master_read_data_valid_sdram_s1_shift_register),
      .cpu_instruction_master_requests_cpu_jtag_debug_module          (cpu_instruction_master_requests_cpu_jtag_debug_module),
      .cpu_jtag_debug_module_address                                  (cpu_jtag_debug_module_address),
      .cpu_jtag_debug_module_begintransfer                            (cpu_jtag_debug_module_begintransfer),
      .cpu_jtag_debug_module_byteenable                               (cpu_jtag_debug_module_byteenable),
      .cpu_jtag_debug_module_chipselect                               (cpu_jtag_debug_module_chipselect),
      .cpu_jtag_debug_module_debugaccess                              (cpu_jtag_debug_module_debugaccess),
      .cpu_jtag_debug_module_readdata                                 (cpu_jtag_debug_module_readdata),
      .cpu_jtag_debug_module_readdata_from_sa                         (cpu_jtag_debug_module_readdata_from_sa),
      .cpu_jtag_debug_module_reset_n                                  (cpu_jtag_debug_module_reset_n),
      .cpu_jtag_debug_module_resetrequest                             (cpu_jtag_debug_module_resetrequest),
      .cpu_jtag_debug_module_resetrequest_from_sa                     (cpu_jtag_debug_module_resetrequest_from_sa),
      .cpu_jtag_debug_module_write                                    (cpu_jtag_debug_module_write),
      .cpu_jtag_debug_module_writedata                                (cpu_jtag_debug_module_writedata),
      .d1_cpu_jtag_debug_module_end_xfer                              (d1_cpu_jtag_debug_module_end_xfer),
      .reset_n                                                        (clk_reset_n)
    );

  cpu_data_master_arbitrator the_cpu_data_master
    (
      .PIO_LCD_B_s1_readdata_from_sa                                 (PIO_LCD_B_s1_readdata_from_sa),
      .PIO_LCD_CLK_s1_readdata_from_sa                               (PIO_LCD_CLK_s1_readdata_from_sa),
      .PIO_LCD_CTRL_s1_readdata_from_sa                              (PIO_LCD_CTRL_s1_readdata_from_sa),
      .PIO_LCD_G_s1_readdata_from_sa                                 (PIO_LCD_G_s1_readdata_from_sa),
      .PIO_LCD_PWM_s1_readdata_from_sa                               (PIO_LCD_PWM_s1_readdata_from_sa),
      .PIO_LCD_R_s1_readdata_from_sa                                 (PIO_LCD_R_s1_readdata_from_sa),
      .PIO_LED_s1_readdata_from_sa                                   (PIO_LED_s1_readdata_from_sa),
      .RS232_s1_irq_from_sa                                          (RS232_s1_irq_from_sa),
      .RS232_s1_readdata_from_sa                                     (RS232_s1_readdata_from_sa),
      .clk                                                           (clk),
      .cpu_data_master_address                                       (cpu_data_master_address),
      .cpu_data_master_address_to_slave                              (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable_sdram_s1                           (cpu_data_master_byteenable_sdram_s1),
      .cpu_data_master_dbs_address                                   (cpu_data_master_dbs_address),
      .cpu_data_master_dbs_write_16                                  (cpu_data_master_dbs_write_16),
      .cpu_data_master_granted_PIO_LCD_B_s1                          (cpu_data_master_granted_PIO_LCD_B_s1),
      .cpu_data_master_granted_PIO_LCD_CLK_s1                        (cpu_data_master_granted_PIO_LCD_CLK_s1),
      .cpu_data_master_granted_PIO_LCD_CTRL_s1                       (cpu_data_master_granted_PIO_LCD_CTRL_s1),
      .cpu_data_master_granted_PIO_LCD_G_s1                          (cpu_data_master_granted_PIO_LCD_G_s1),
      .cpu_data_master_granted_PIO_LCD_PWM_s1                        (cpu_data_master_granted_PIO_LCD_PWM_s1),
      .cpu_data_master_granted_PIO_LCD_R_s1                          (cpu_data_master_granted_PIO_LCD_R_s1),
      .cpu_data_master_granted_PIO_LED_s1                            (cpu_data_master_granted_PIO_LED_s1),
      .cpu_data_master_granted_RS232_s1                              (cpu_data_master_granted_RS232_s1),
      .cpu_data_master_granted_cpu_jtag_debug_module                 (cpu_data_master_granted_cpu_jtag_debug_module),
      .cpu_data_master_granted_epcs_epcs_control_port                (cpu_data_master_granted_epcs_epcs_control_port),
      .cpu_data_master_granted_jtag_uart_avalon_jtag_slave           (cpu_data_master_granted_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_granted_sdram_s1                              (cpu_data_master_granted_sdram_s1),
      .cpu_data_master_granted_sysid_control_slave                   (cpu_data_master_granted_sysid_control_slave),
      .cpu_data_master_irq                                           (cpu_data_master_irq),
      .cpu_data_master_no_byte_enables_and_last_term                 (cpu_data_master_no_byte_enables_and_last_term),
      .cpu_data_master_qualified_request_PIO_LCD_B_s1                (cpu_data_master_qualified_request_PIO_LCD_B_s1),
      .cpu_data_master_qualified_request_PIO_LCD_CLK_s1              (cpu_data_master_qualified_request_PIO_LCD_CLK_s1),
      .cpu_data_master_qualified_request_PIO_LCD_CTRL_s1             (cpu_data_master_qualified_request_PIO_LCD_CTRL_s1),
      .cpu_data_master_qualified_request_PIO_LCD_G_s1                (cpu_data_master_qualified_request_PIO_LCD_G_s1),
      .cpu_data_master_qualified_request_PIO_LCD_PWM_s1              (cpu_data_master_qualified_request_PIO_LCD_PWM_s1),
      .cpu_data_master_qualified_request_PIO_LCD_R_s1                (cpu_data_master_qualified_request_PIO_LCD_R_s1),
      .cpu_data_master_qualified_request_PIO_LED_s1                  (cpu_data_master_qualified_request_PIO_LED_s1),
      .cpu_data_master_qualified_request_RS232_s1                    (cpu_data_master_qualified_request_RS232_s1),
      .cpu_data_master_qualified_request_cpu_jtag_debug_module       (cpu_data_master_qualified_request_cpu_jtag_debug_module),
      .cpu_data_master_qualified_request_epcs_epcs_control_port      (cpu_data_master_qualified_request_epcs_epcs_control_port),
      .cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave (cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_qualified_request_sdram_s1                    (cpu_data_master_qualified_request_sdram_s1),
      .cpu_data_master_qualified_request_sysid_control_slave         (cpu_data_master_qualified_request_sysid_control_slave),
      .cpu_data_master_read                                          (cpu_data_master_read),
      .cpu_data_master_read_data_valid_PIO_LCD_B_s1                  (cpu_data_master_read_data_valid_PIO_LCD_B_s1),
      .cpu_data_master_read_data_valid_PIO_LCD_CLK_s1                (cpu_data_master_read_data_valid_PIO_LCD_CLK_s1),
      .cpu_data_master_read_data_valid_PIO_LCD_CTRL_s1               (cpu_data_master_read_data_valid_PIO_LCD_CTRL_s1),
      .cpu_data_master_read_data_valid_PIO_LCD_G_s1                  (cpu_data_master_read_data_valid_PIO_LCD_G_s1),
      .cpu_data_master_read_data_valid_PIO_LCD_PWM_s1                (cpu_data_master_read_data_valid_PIO_LCD_PWM_s1),
      .cpu_data_master_read_data_valid_PIO_LCD_R_s1                  (cpu_data_master_read_data_valid_PIO_LCD_R_s1),
      .cpu_data_master_read_data_valid_PIO_LED_s1                    (cpu_data_master_read_data_valid_PIO_LED_s1),
      .cpu_data_master_read_data_valid_RS232_s1                      (cpu_data_master_read_data_valid_RS232_s1),
      .cpu_data_master_read_data_valid_cpu_jtag_debug_module         (cpu_data_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_data_master_read_data_valid_epcs_epcs_control_port        (cpu_data_master_read_data_valid_epcs_epcs_control_port),
      .cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave   (cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_read_data_valid_sdram_s1                      (cpu_data_master_read_data_valid_sdram_s1),
      .cpu_data_master_read_data_valid_sdram_s1_shift_register       (cpu_data_master_read_data_valid_sdram_s1_shift_register),
      .cpu_data_master_read_data_valid_sysid_control_slave           (cpu_data_master_read_data_valid_sysid_control_slave),
      .cpu_data_master_readdata                                      (cpu_data_master_readdata),
      .cpu_data_master_requests_PIO_LCD_B_s1                         (cpu_data_master_requests_PIO_LCD_B_s1),
      .cpu_data_master_requests_PIO_LCD_CLK_s1                       (cpu_data_master_requests_PIO_LCD_CLK_s1),
      .cpu_data_master_requests_PIO_LCD_CTRL_s1                      (cpu_data_master_requests_PIO_LCD_CTRL_s1),
      .cpu_data_master_requests_PIO_LCD_G_s1                         (cpu_data_master_requests_PIO_LCD_G_s1),
      .cpu_data_master_requests_PIO_LCD_PWM_s1                       (cpu_data_master_requests_PIO_LCD_PWM_s1),
      .cpu_data_master_requests_PIO_LCD_R_s1                         (cpu_data_master_requests_PIO_LCD_R_s1),
      .cpu_data_master_requests_PIO_LED_s1                           (cpu_data_master_requests_PIO_LED_s1),
      .cpu_data_master_requests_RS232_s1                             (cpu_data_master_requests_RS232_s1),
      .cpu_data_master_requests_cpu_jtag_debug_module                (cpu_data_master_requests_cpu_jtag_debug_module),
      .cpu_data_master_requests_epcs_epcs_control_port               (cpu_data_master_requests_epcs_epcs_control_port),
      .cpu_data_master_requests_jtag_uart_avalon_jtag_slave          (cpu_data_master_requests_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_requests_sdram_s1                             (cpu_data_master_requests_sdram_s1),
      .cpu_data_master_requests_sysid_control_slave                  (cpu_data_master_requests_sysid_control_slave),
      .cpu_data_master_waitrequest                                   (cpu_data_master_waitrequest),
      .cpu_data_master_write                                         (cpu_data_master_write),
      .cpu_data_master_writedata                                     (cpu_data_master_writedata),
      .cpu_jtag_debug_module_readdata_from_sa                        (cpu_jtag_debug_module_readdata_from_sa),
      .d1_PIO_LCD_B_s1_end_xfer                                      (d1_PIO_LCD_B_s1_end_xfer),
      .d1_PIO_LCD_CLK_s1_end_xfer                                    (d1_PIO_LCD_CLK_s1_end_xfer),
      .d1_PIO_LCD_CTRL_s1_end_xfer                                   (d1_PIO_LCD_CTRL_s1_end_xfer),
      .d1_PIO_LCD_G_s1_end_xfer                                      (d1_PIO_LCD_G_s1_end_xfer),
      .d1_PIO_LCD_PWM_s1_end_xfer                                    (d1_PIO_LCD_PWM_s1_end_xfer),
      .d1_PIO_LCD_R_s1_end_xfer                                      (d1_PIO_LCD_R_s1_end_xfer),
      .d1_PIO_LED_s1_end_xfer                                        (d1_PIO_LED_s1_end_xfer),
      .d1_RS232_s1_end_xfer                                          (d1_RS232_s1_end_xfer),
      .d1_cpu_jtag_debug_module_end_xfer                             (d1_cpu_jtag_debug_module_end_xfer),
      .d1_epcs_epcs_control_port_end_xfer                            (d1_epcs_epcs_control_port_end_xfer),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                       (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .d1_sdram_s1_end_xfer                                          (d1_sdram_s1_end_xfer),
      .d1_sysid_control_slave_end_xfer                               (d1_sysid_control_slave_end_xfer),
      .epcs_epcs_control_port_irq_from_sa                            (epcs_epcs_control_port_irq_from_sa),
      .epcs_epcs_control_port_readdata_from_sa                       (epcs_epcs_control_port_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                       (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                  (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa               (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .reset_n                                                       (clk_reset_n),
      .sdram_s1_readdata_from_sa                                     (sdram_s1_readdata_from_sa),
      .sdram_s1_waitrequest_from_sa                                  (sdram_s1_waitrequest_from_sa),
      .sysid_control_slave_readdata_from_sa                          (sysid_control_slave_readdata_from_sa)
    );

  cpu_instruction_master_arbitrator the_cpu_instruction_master
    (
      .clk                                                             (clk),
      .cpu_instruction_master_address                                  (cpu_instruction_master_address),
      .cpu_instruction_master_address_to_slave                         (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_dbs_address                              (cpu_instruction_master_dbs_address),
      .cpu_instruction_master_granted_cpu_jtag_debug_module            (cpu_instruction_master_granted_cpu_jtag_debug_module),
      .cpu_instruction_master_granted_epcs_epcs_control_port           (cpu_instruction_master_granted_epcs_epcs_control_port),
      .cpu_instruction_master_granted_sdram_s1                         (cpu_instruction_master_granted_sdram_s1),
      .cpu_instruction_master_latency_counter                          (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_cpu_jtag_debug_module  (cpu_instruction_master_qualified_request_cpu_jtag_debug_module),
      .cpu_instruction_master_qualified_request_epcs_epcs_control_port (cpu_instruction_master_qualified_request_epcs_epcs_control_port),
      .cpu_instruction_master_qualified_request_sdram_s1               (cpu_instruction_master_qualified_request_sdram_s1),
      .cpu_instruction_master_read                                     (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_cpu_jtag_debug_module    (cpu_instruction_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_instruction_master_read_data_valid_epcs_epcs_control_port   (cpu_instruction_master_read_data_valid_epcs_epcs_control_port),
      .cpu_instruction_master_read_data_valid_sdram_s1                 (cpu_instruction_master_read_data_valid_sdram_s1),
      .cpu_instruction_master_read_data_valid_sdram_s1_shift_register  (cpu_instruction_master_read_data_valid_sdram_s1_shift_register),
      .cpu_instruction_master_readdata                                 (cpu_instruction_master_readdata),
      .cpu_instruction_master_readdatavalid                            (cpu_instruction_master_readdatavalid),
      .cpu_instruction_master_requests_cpu_jtag_debug_module           (cpu_instruction_master_requests_cpu_jtag_debug_module),
      .cpu_instruction_master_requests_epcs_epcs_control_port          (cpu_instruction_master_requests_epcs_epcs_control_port),
      .cpu_instruction_master_requests_sdram_s1                        (cpu_instruction_master_requests_sdram_s1),
      .cpu_instruction_master_waitrequest                              (cpu_instruction_master_waitrequest),
      .cpu_jtag_debug_module_readdata_from_sa                          (cpu_jtag_debug_module_readdata_from_sa),
      .d1_cpu_jtag_debug_module_end_xfer                               (d1_cpu_jtag_debug_module_end_xfer),
      .d1_epcs_epcs_control_port_end_xfer                              (d1_epcs_epcs_control_port_end_xfer),
      .d1_sdram_s1_end_xfer                                            (d1_sdram_s1_end_xfer),
      .epcs_epcs_control_port_readdata_from_sa                         (epcs_epcs_control_port_readdata_from_sa),
      .reset_n                                                         (clk_reset_n),
      .sdram_s1_readdata_from_sa                                       (sdram_s1_readdata_from_sa),
      .sdram_s1_waitrequest_from_sa                                    (sdram_s1_waitrequest_from_sa)
    );

  cpu the_cpu
    (
      .clk                                   (clk),
      .d_address                             (cpu_data_master_address),
      .d_byteenable                          (cpu_data_master_byteenable),
      .d_irq                                 (cpu_data_master_irq),
      .d_read                                (cpu_data_master_read),
      .d_readdata                            (cpu_data_master_readdata),
      .d_waitrequest                         (cpu_data_master_waitrequest),
      .d_write                               (cpu_data_master_write),
      .d_writedata                           (cpu_data_master_writedata),
      .i_address                             (cpu_instruction_master_address),
      .i_read                                (cpu_instruction_master_read),
      .i_readdata                            (cpu_instruction_master_readdata),
      .i_readdatavalid                       (cpu_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_instruction_master_waitrequest),
      .jtag_debug_module_address             (cpu_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_jtag_debug_module_byteenable),
      .jtag_debug_module_debugaccess         (cpu_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_jtag_debug_module_readdata),
      .jtag_debug_module_resetrequest        (cpu_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_jtag_debug_module_writedata),
      .reset_n                               (cpu_jtag_debug_module_reset_n)
    );

  epcs_epcs_control_port_arbitrator the_epcs_epcs_control_port
    (
      .clk                                                             (clk),
      .cpu_data_master_address_to_slave                                (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_epcs_epcs_control_port                  (cpu_data_master_granted_epcs_epcs_control_port),
      .cpu_data_master_qualified_request_epcs_epcs_control_port        (cpu_data_master_qualified_request_epcs_epcs_control_port),
      .cpu_data_master_read                                            (cpu_data_master_read),
      .cpu_data_master_read_data_valid_epcs_epcs_control_port          (cpu_data_master_read_data_valid_epcs_epcs_control_port),
      .cpu_data_master_requests_epcs_epcs_control_port                 (cpu_data_master_requests_epcs_epcs_control_port),
      .cpu_data_master_write                                           (cpu_data_master_write),
      .cpu_data_master_writedata                                       (cpu_data_master_writedata),
      .cpu_instruction_master_address_to_slave                         (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_epcs_epcs_control_port           (cpu_instruction_master_granted_epcs_epcs_control_port),
      .cpu_instruction_master_latency_counter                          (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_epcs_epcs_control_port (cpu_instruction_master_qualified_request_epcs_epcs_control_port),
      .cpu_instruction_master_read                                     (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_epcs_epcs_control_port   (cpu_instruction_master_read_data_valid_epcs_epcs_control_port),
      .cpu_instruction_master_read_data_valid_sdram_s1_shift_register  (cpu_instruction_master_read_data_valid_sdram_s1_shift_register),
      .cpu_instruction_master_requests_epcs_epcs_control_port          (cpu_instruction_master_requests_epcs_epcs_control_port),
      .d1_epcs_epcs_control_port_end_xfer                              (d1_epcs_epcs_control_port_end_xfer),
      .epcs_epcs_control_port_address                                  (epcs_epcs_control_port_address),
      .epcs_epcs_control_port_chipselect                               (epcs_epcs_control_port_chipselect),
      .epcs_epcs_control_port_dataavailable                            (epcs_epcs_control_port_dataavailable),
      .epcs_epcs_control_port_dataavailable_from_sa                    (epcs_epcs_control_port_dataavailable_from_sa),
      .epcs_epcs_control_port_endofpacket                              (epcs_epcs_control_port_endofpacket),
      .epcs_epcs_control_port_endofpacket_from_sa                      (epcs_epcs_control_port_endofpacket_from_sa),
      .epcs_epcs_control_port_irq                                      (epcs_epcs_control_port_irq),
      .epcs_epcs_control_port_irq_from_sa                              (epcs_epcs_control_port_irq_from_sa),
      .epcs_epcs_control_port_read_n                                   (epcs_epcs_control_port_read_n),
      .epcs_epcs_control_port_readdata                                 (epcs_epcs_control_port_readdata),
      .epcs_epcs_control_port_readdata_from_sa                         (epcs_epcs_control_port_readdata_from_sa),
      .epcs_epcs_control_port_readyfordata                             (epcs_epcs_control_port_readyfordata),
      .epcs_epcs_control_port_readyfordata_from_sa                     (epcs_epcs_control_port_readyfordata_from_sa),
      .epcs_epcs_control_port_reset_n                                  (epcs_epcs_control_port_reset_n),
      .epcs_epcs_control_port_write_n                                  (epcs_epcs_control_port_write_n),
      .epcs_epcs_control_port_writedata                                (epcs_epcs_control_port_writedata),
      .reset_n                                                         (clk_reset_n)
    );

  epcs the_epcs
    (
      .address       (epcs_epcs_control_port_address),
      .chipselect    (epcs_epcs_control_port_chipselect),
      .clk           (clk),
      .data0         (data0_to_the_epcs),
      .dataavailable (epcs_epcs_control_port_dataavailable),
      .dclk          (dclk_from_the_epcs),
      .endofpacket   (epcs_epcs_control_port_endofpacket),
      .irq           (epcs_epcs_control_port_irq),
      .read_n        (epcs_epcs_control_port_read_n),
      .readdata      (epcs_epcs_control_port_readdata),
      .readyfordata  (epcs_epcs_control_port_readyfordata),
      .reset_n       (epcs_epcs_control_port_reset_n),
      .sce           (sce_from_the_epcs),
      .sdo           (sdo_from_the_epcs),
      .write_n       (epcs_epcs_control_port_write_n),
      .writedata     (epcs_epcs_control_port_writedata)
    );

  jtag_uart_avalon_jtag_slave_arbitrator the_jtag_uart_avalon_jtag_slave
    (
      .clk                                                           (clk),
      .cpu_data_master_address_to_slave                              (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_jtag_uart_avalon_jtag_slave           (cpu_data_master_granted_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave (cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_read                                          (cpu_data_master_read),
      .cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave   (cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_requests_jtag_uart_avalon_jtag_slave          (cpu_data_master_requests_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_waitrequest                                   (cpu_data_master_waitrequest),
      .cpu_data_master_write                                         (cpu_data_master_write),
      .cpu_data_master_writedata                                     (cpu_data_master_writedata),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                       (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .jtag_uart_avalon_jtag_slave_address                           (jtag_uart_avalon_jtag_slave_address),
      .jtag_uart_avalon_jtag_slave_chipselect                        (jtag_uart_avalon_jtag_slave_chipselect),
      .jtag_uart_avalon_jtag_slave_dataavailable                     (jtag_uart_avalon_jtag_slave_dataavailable),
      .jtag_uart_avalon_jtag_slave_dataavailable_from_sa             (jtag_uart_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_avalon_jtag_slave_irq                               (jtag_uart_avalon_jtag_slave_irq),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                       (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_read_n                            (jtag_uart_avalon_jtag_slave_read_n),
      .jtag_uart_avalon_jtag_slave_readdata                          (jtag_uart_avalon_jtag_slave_readdata),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                  (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_readyfordata                      (jtag_uart_avalon_jtag_slave_readyfordata),
      .jtag_uart_avalon_jtag_slave_readyfordata_from_sa              (jtag_uart_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_avalon_jtag_slave_reset_n                           (jtag_uart_avalon_jtag_slave_reset_n),
      .jtag_uart_avalon_jtag_slave_waitrequest                       (jtag_uart_avalon_jtag_slave_waitrequest),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa               (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_avalon_jtag_slave_write_n                           (jtag_uart_avalon_jtag_slave_write_n),
      .jtag_uart_avalon_jtag_slave_writedata                         (jtag_uart_avalon_jtag_slave_writedata),
      .reset_n                                                       (clk_reset_n)
    );

  jtag_uart the_jtag_uart
    (
      .av_address     (jtag_uart_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_avalon_jtag_slave_writedata),
      .clk            (clk),
      .dataavailable  (jtag_uart_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_avalon_jtag_slave_reset_n)
    );

  sdram_s1_arbitrator the_sdram_s1
    (
      .clk                                                            (clk),
      .cpu_data_master_address_to_slave                               (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                     (cpu_data_master_byteenable),
      .cpu_data_master_byteenable_sdram_s1                            (cpu_data_master_byteenable_sdram_s1),
      .cpu_data_master_dbs_address                                    (cpu_data_master_dbs_address),
      .cpu_data_master_dbs_write_16                                   (cpu_data_master_dbs_write_16),
      .cpu_data_master_granted_sdram_s1                               (cpu_data_master_granted_sdram_s1),
      .cpu_data_master_no_byte_enables_and_last_term                  (cpu_data_master_no_byte_enables_and_last_term),
      .cpu_data_master_qualified_request_sdram_s1                     (cpu_data_master_qualified_request_sdram_s1),
      .cpu_data_master_read                                           (cpu_data_master_read),
      .cpu_data_master_read_data_valid_sdram_s1                       (cpu_data_master_read_data_valid_sdram_s1),
      .cpu_data_master_read_data_valid_sdram_s1_shift_register        (cpu_data_master_read_data_valid_sdram_s1_shift_register),
      .cpu_data_master_requests_sdram_s1                              (cpu_data_master_requests_sdram_s1),
      .cpu_data_master_waitrequest                                    (cpu_data_master_waitrequest),
      .cpu_data_master_write                                          (cpu_data_master_write),
      .cpu_instruction_master_address_to_slave                        (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_dbs_address                             (cpu_instruction_master_dbs_address),
      .cpu_instruction_master_granted_sdram_s1                        (cpu_instruction_master_granted_sdram_s1),
      .cpu_instruction_master_latency_counter                         (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_sdram_s1              (cpu_instruction_master_qualified_request_sdram_s1),
      .cpu_instruction_master_read                                    (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_sdram_s1                (cpu_instruction_master_read_data_valid_sdram_s1),
      .cpu_instruction_master_read_data_valid_sdram_s1_shift_register (cpu_instruction_master_read_data_valid_sdram_s1_shift_register),
      .cpu_instruction_master_requests_sdram_s1                       (cpu_instruction_master_requests_sdram_s1),
      .d1_sdram_s1_end_xfer                                           (d1_sdram_s1_end_xfer),
      .reset_n                                                        (clk_reset_n),
      .sdram_s1_address                                               (sdram_s1_address),
      .sdram_s1_byteenable_n                                          (sdram_s1_byteenable_n),
      .sdram_s1_chipselect                                            (sdram_s1_chipselect),
      .sdram_s1_read_n                                                (sdram_s1_read_n),
      .sdram_s1_readdata                                              (sdram_s1_readdata),
      .sdram_s1_readdata_from_sa                                      (sdram_s1_readdata_from_sa),
      .sdram_s1_readdatavalid                                         (sdram_s1_readdatavalid),
      .sdram_s1_reset_n                                               (sdram_s1_reset_n),
      .sdram_s1_waitrequest                                           (sdram_s1_waitrequest),
      .sdram_s1_waitrequest_from_sa                                   (sdram_s1_waitrequest_from_sa),
      .sdram_s1_write_n                                               (sdram_s1_write_n),
      .sdram_s1_writedata                                             (sdram_s1_writedata)
    );

  sdram the_sdram
    (
      .az_addr        (sdram_s1_address),
      .az_be_n        (sdram_s1_byteenable_n),
      .az_cs          (sdram_s1_chipselect),
      .az_data        (sdram_s1_writedata),
      .az_rd_n        (sdram_s1_read_n),
      .az_wr_n        (sdram_s1_write_n),
      .clk            (clk),
      .reset_n        (sdram_s1_reset_n),
      .za_data        (sdram_s1_readdata),
      .za_valid       (sdram_s1_readdatavalid),
      .za_waitrequest (sdram_s1_waitrequest),
      .zs_addr        (zs_addr_from_the_sdram),
      .zs_ba          (zs_ba_from_the_sdram),
      .zs_cas_n       (zs_cas_n_from_the_sdram),
      .zs_cke         (zs_cke_from_the_sdram),
      .zs_cs_n        (zs_cs_n_from_the_sdram),
      .zs_dq          (zs_dq_to_and_from_the_sdram),
      .zs_dqm         (zs_dqm_from_the_sdram),
      .zs_ras_n       (zs_ras_n_from_the_sdram),
      .zs_we_n        (zs_we_n_from_the_sdram)
    );

  sysid_control_slave_arbitrator the_sysid_control_slave
    (
      .clk                                                   (clk),
      .cpu_data_master_address_to_slave                      (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_sysid_control_slave           (cpu_data_master_granted_sysid_control_slave),
      .cpu_data_master_qualified_request_sysid_control_slave (cpu_data_master_qualified_request_sysid_control_slave),
      .cpu_data_master_read                                  (cpu_data_master_read),
      .cpu_data_master_read_data_valid_sysid_control_slave   (cpu_data_master_read_data_valid_sysid_control_slave),
      .cpu_data_master_requests_sysid_control_slave          (cpu_data_master_requests_sysid_control_slave),
      .cpu_data_master_write                                 (cpu_data_master_write),
      .d1_sysid_control_slave_end_xfer                       (d1_sysid_control_slave_end_xfer),
      .reset_n                                               (clk_reset_n),
      .sysid_control_slave_address                           (sysid_control_slave_address),
      .sysid_control_slave_readdata                          (sysid_control_slave_readdata),
      .sysid_control_slave_readdata_from_sa                  (sysid_control_slave_readdata_from_sa),
      .sysid_control_slave_reset_n                           (sysid_control_slave_reset_n)
    );

  sysid the_sysid
    (
      .address  (sysid_control_slave_address),
      .clock    (sysid_control_slave_clock),
      .readdata (sysid_control_slave_readdata),
      .reset_n  (sysid_control_slave_reset_n)
    );

  //reset is asserted asynchronously and deasserted synchronously
  kernel_reset_clk_domain_synch_module kernel_reset_clk_domain_synch
    (
      .clk      (clk),
      .data_in  (1'b1),
      .data_out (clk_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset sources mux, which is an e_mux
  assign reset_n_sources = ~(~reset_n |
    0 |
    cpu_jtag_debug_module_resetrequest_from_sa |
    cpu_jtag_debug_module_resetrequest_from_sa);

  //sysid_control_slave_clock of type clock does not connect to anything so wire it to default (0)
  assign sysid_control_slave_clock = 0;


endmodule


//synthesis translate_off



// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE

// AND HERE WILL BE PRESERVED </ALTERA_NOTE>


// If user logic components use Altsync_Ram with convert_hex2ver.dll,
// set USE_convert_hex2ver in the user comments section above

// `ifdef USE_convert_hex2ver
// `else
// `define NO_PLI 1
// `endif

`include "c:/altera/11.0/quartus/eda/sim_lib/altera_mf.v"
`include "c:/altera/11.0/quartus/eda/sim_lib/220model.v"
`include "c:/altera/11.0/quartus/eda/sim_lib/sgate.v"
`include "PIO_LCD_G.v"
`include "PIO_LCD_PWM.v"
`include "cpu_test_bench.v"
`include "cpu_mult_cell.v"
`include "cpu_oci_test_bench.v"
`include "cpu_jtag_debug_module_tck.v"
`include "cpu_jtag_debug_module_sysclk.v"
`include "cpu_jtag_debug_module_wrapper.v"
`include "cpu.v"
`include "sdram.v"
`include "sysid.v"
`include "PIO_LCD_R.v"
`include "PIO_LED.v"
`include "epcs.v"
`include "jtag_uart.v"
`include "PIO_LCD_CTRL.v"
`include "PIO_LCD_CLK.v"
`include "PIO_LCD_B.v"
`include "RS232.v"

`timescale 1ns / 1ps

module test_bench 
;


  wire             RS232_s1_dataavailable_from_sa;
  wire             RS232_s1_readyfordata_from_sa;
  reg              clk;
  wire             data0_to_the_epcs;
  wire             dclk_from_the_epcs;
  wire             epcs_epcs_control_port_dataavailable_from_sa;
  wire             epcs_epcs_control_port_endofpacket_from_sa;
  wire             epcs_epcs_control_port_readyfordata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire    [  5: 0] out_port_from_the_PIO_LCD_B;
  wire             out_port_from_the_PIO_LCD_CLK;
  wire    [  7: 0] out_port_from_the_PIO_LCD_CTRL;
  wire    [  5: 0] out_port_from_the_PIO_LCD_G;
  wire             out_port_from_the_PIO_LCD_PWM;
  wire    [  5: 0] out_port_from_the_PIO_LCD_R;
  wire    [  3: 0] out_port_from_the_PIO_LED;
  reg              reset_n;
  wire             rxd_to_the_RS232;
  wire             sce_from_the_epcs;
  wire             sdo_from_the_epcs;
  wire             sysid_control_slave_clock;
  wire             txd_from_the_RS232;
  wire    [ 12: 0] zs_addr_from_the_sdram;
  wire    [  1: 0] zs_ba_from_the_sdram;
  wire             zs_cas_n_from_the_sdram;
  wire             zs_cke_from_the_sdram;
  wire             zs_cs_n_from_the_sdram;
  wire    [ 15: 0] zs_dq_to_and_from_the_sdram;
  wire    [  1: 0] zs_dqm_from_the_sdram;
  wire             zs_ras_n_from_the_sdram;
  wire             zs_we_n_from_the_sdram;


// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
//  add your signals and additional architecture here
// AND HERE WILL BE PRESERVED </ALTERA_NOTE>

  //Set us up the Dut
  kernel DUT
    (
      .clk                            (clk),
      .data0_to_the_epcs              (data0_to_the_epcs),
      .dclk_from_the_epcs             (dclk_from_the_epcs),
      .out_port_from_the_PIO_LCD_B    (out_port_from_the_PIO_LCD_B),
      .out_port_from_the_PIO_LCD_CLK  (out_port_from_the_PIO_LCD_CLK),
      .out_port_from_the_PIO_LCD_CTRL (out_port_from_the_PIO_LCD_CTRL),
      .out_port_from_the_PIO_LCD_G    (out_port_from_the_PIO_LCD_G),
      .out_port_from_the_PIO_LCD_PWM  (out_port_from_the_PIO_LCD_PWM),
      .out_port_from_the_PIO_LCD_R    (out_port_from_the_PIO_LCD_R),
      .out_port_from_the_PIO_LED      (out_port_from_the_PIO_LED),
      .reset_n                        (reset_n),
      .rxd_to_the_RS232               (rxd_to_the_RS232),
      .sce_from_the_epcs              (sce_from_the_epcs),
      .sdo_from_the_epcs              (sdo_from_the_epcs),
      .txd_from_the_RS232             (txd_from_the_RS232),
      .zs_addr_from_the_sdram         (zs_addr_from_the_sdram),
      .zs_ba_from_the_sdram           (zs_ba_from_the_sdram),
      .zs_cas_n_from_the_sdram        (zs_cas_n_from_the_sdram),
      .zs_cke_from_the_sdram          (zs_cke_from_the_sdram),
      .zs_cs_n_from_the_sdram         (zs_cs_n_from_the_sdram),
      .zs_dq_to_and_from_the_sdram    (zs_dq_to_and_from_the_sdram),
      .zs_dqm_from_the_sdram          (zs_dqm_from_the_sdram),
      .zs_ras_n_from_the_sdram        (zs_ras_n_from_the_sdram),
      .zs_we_n_from_the_sdram         (zs_we_n_from_the_sdram)
    );

  initial
    clk = 1'b0;
  always
    #5 clk <= ~clk;
  
  initial 
    begin
      reset_n <= 0;
      #100 reset_n <= 1;
    end

endmodule


//synthesis translate_on