module main;
initial 
begin 
	$display("helloworld");
	$finish;
end 
endmodule
