module counter;
initial 
begin 
	$display("helloworld");
	$finish;
end 
endmodule
